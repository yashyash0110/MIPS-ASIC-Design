VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cpu
  CLASS BLOCK ;
  FOREIGN cpu ;
  ORIGIN 0.000 0.000 ;
  SIZE 125.000 BY 135.720 ;
  PIN MEM_WRITE[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END MEM_WRITE[0]
  PIN MEM_WRITE[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END MEM_WRITE[10]
  PIN MEM_WRITE[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END MEM_WRITE[11]
  PIN MEM_WRITE[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 131.720 55.110 135.720 ;
    END
  END MEM_WRITE[12]
  PIN MEM_WRITE[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END MEM_WRITE[13]
  PIN MEM_WRITE[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 131.720 42.230 135.720 ;
    END
  END MEM_WRITE[14]
  PIN MEM_WRITE[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 131.720 39.010 135.720 ;
    END
  END MEM_WRITE[15]
  PIN MEM_WRITE[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 67.710 131.720 67.990 135.720 ;
    END
  END MEM_WRITE[16]
  PIN MEM_WRITE[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 70.930 131.720 71.210 135.720 ;
    END
  END MEM_WRITE[17]
  PIN MEM_WRITE[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 121.000 68.040 125.000 68.640 ;
    END
  END MEM_WRITE[18]
  PIN MEM_WRITE[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 131.720 74.430 135.720 ;
    END
  END MEM_WRITE[19]
  PIN MEM_WRITE[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 121.000 61.240 125.000 61.840 ;
    END
  END MEM_WRITE[1]
  PIN MEM_WRITE[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 121.000 95.240 125.000 95.840 ;
    END
  END MEM_WRITE[20]
  PIN MEM_WRITE[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 121.000 91.840 125.000 92.440 ;
    END
  END MEM_WRITE[21]
  PIN MEM_WRITE[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 121.000 81.640 125.000 82.240 ;
    END
  END MEM_WRITE[22]
  PIN MEM_WRITE[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 121.000 78.240 125.000 78.840 ;
    END
  END MEM_WRITE[23]
  PIN MEM_WRITE[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 121.000 64.640 125.000 65.240 ;
    END
  END MEM_WRITE[24]
  PIN MEM_WRITE[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 121.000 71.440 125.000 72.040 ;
    END
  END MEM_WRITE[25]
  PIN MEM_WRITE[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 121.000 54.440 125.000 55.040 ;
    END
  END MEM_WRITE[26]
  PIN MEM_WRITE[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 121.000 57.840 125.000 58.440 ;
    END
  END MEM_WRITE[27]
  PIN MEM_WRITE[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 121.000 44.240 125.000 44.840 ;
    END
  END MEM_WRITE[28]
  PIN MEM_WRITE[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 121.000 40.840 125.000 41.440 ;
    END
  END MEM_WRITE[29]
  PIN MEM_WRITE[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END MEM_WRITE[2]
  PIN MEM_WRITE[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END MEM_WRITE[30]
  PIN MEM_WRITE[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END MEM_WRITE[31]
  PIN MEM_WRITE[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END MEM_WRITE[3]
  PIN MEM_WRITE[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END MEM_WRITE[4]
  PIN MEM_WRITE[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END MEM_WRITE[5]
  PIN MEM_WRITE[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END MEM_WRITE[6]
  PIN MEM_WRITE[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END MEM_WRITE[7]
  PIN MEM_WRITE[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END MEM_WRITE[8]
  PIN MEM_WRITE[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END MEM_WRITE[9]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -5.380 -0.020 -3.780 133.300 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 -0.020 130.040 1.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 131.700 130.040 133.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 128.440 -0.020 130.040 133.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 13.220 -0.020 15.220 133.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 43.220 -0.020 45.220 133.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.220 -0.020 75.220 133.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 103.220 -0.020 105.220 133.300 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 18.580 130.040 20.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 48.580 130.040 50.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 78.580 130.040 80.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 108.580 130.040 110.580 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -2.080 3.280 -0.480 130.000 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 3.280 126.740 4.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 128.400 126.740 130.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.140 3.280 126.740 130.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.520 -0.020 11.520 133.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.520 -0.020 41.520 133.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.520 -0.020 71.520 133.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.520 -0.020 101.520 133.300 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 14.880 130.040 16.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 44.880 130.040 46.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 74.880 130.040 76.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 104.880 130.040 106.880 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END rst
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 119.140 122.485 ;
      LAYER met1 ;
        RECT 4.670 10.640 119.140 122.640 ;
      LAYER met2 ;
        RECT 4.690 131.440 38.450 132.330 ;
        RECT 39.290 131.440 41.670 132.330 ;
        RECT 42.510 131.440 54.550 132.330 ;
        RECT 55.390 131.440 67.430 132.330 ;
        RECT 68.270 131.440 70.650 132.330 ;
        RECT 71.490 131.440 73.870 132.330 ;
        RECT 74.710 131.440 117.660 132.330 ;
        RECT 4.690 4.280 117.660 131.440 ;
        RECT 4.690 4.000 35.230 4.280 ;
        RECT 36.070 4.000 38.450 4.280 ;
        RECT 39.290 4.000 51.330 4.280 ;
        RECT 52.170 4.000 54.550 4.280 ;
        RECT 55.390 4.000 60.990 4.280 ;
        RECT 61.830 4.000 64.210 4.280 ;
        RECT 65.050 4.000 67.430 4.280 ;
        RECT 68.270 4.000 86.750 4.280 ;
        RECT 87.590 4.000 89.970 4.280 ;
        RECT 90.810 4.000 117.660 4.280 ;
      LAYER met3 ;
        RECT 4.000 99.640 121.000 122.565 ;
        RECT 4.400 98.240 121.000 99.640 ;
        RECT 4.000 96.240 121.000 98.240 ;
        RECT 4.000 94.840 120.600 96.240 ;
        RECT 4.000 92.840 121.000 94.840 ;
        RECT 4.000 91.440 120.600 92.840 ;
        RECT 4.000 86.040 121.000 91.440 ;
        RECT 4.400 84.640 121.000 86.040 ;
        RECT 4.000 82.640 121.000 84.640 ;
        RECT 4.000 81.240 120.600 82.640 ;
        RECT 4.000 79.240 121.000 81.240 ;
        RECT 4.400 77.840 120.600 79.240 ;
        RECT 4.000 72.440 121.000 77.840 ;
        RECT 4.000 71.040 120.600 72.440 ;
        RECT 4.000 69.040 121.000 71.040 ;
        RECT 4.400 67.640 120.600 69.040 ;
        RECT 4.000 65.640 121.000 67.640 ;
        RECT 4.400 64.240 120.600 65.640 ;
        RECT 4.000 62.240 121.000 64.240 ;
        RECT 4.400 60.840 120.600 62.240 ;
        RECT 4.000 58.840 121.000 60.840 ;
        RECT 4.000 57.440 120.600 58.840 ;
        RECT 4.000 55.440 121.000 57.440 ;
        RECT 4.400 54.040 120.600 55.440 ;
        RECT 4.000 45.240 121.000 54.040 ;
        RECT 4.000 43.840 120.600 45.240 ;
        RECT 4.000 41.840 121.000 43.840 ;
        RECT 4.000 40.440 120.600 41.840 ;
        RECT 4.000 10.715 121.000 40.440 ;
      LAYER met4 ;
        RECT 47.215 53.215 47.545 63.745 ;
  END
END cpu
END LIBRARY

