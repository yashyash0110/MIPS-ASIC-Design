magic
tech sky130A
magscale 1 2
timestamp 1710937663
<< viali >>
rect 8033 24225 8067 24259
rect 9321 24225 9355 24259
rect 11897 24225 11931 24259
rect 14289 24225 14323 24259
rect 15577 24225 15611 24259
rect 7849 24157 7883 24191
rect 9045 24157 9079 24191
rect 11621 24157 11655 24191
rect 14105 24157 14139 24191
rect 14657 24157 14691 24191
rect 14933 24157 14967 24191
rect 15301 24157 15335 24191
rect 11253 22593 11287 22627
rect 11069 22389 11103 22423
rect 9873 22117 9907 22151
rect 9689 22049 9723 22083
rect 8493 21981 8527 22015
rect 8769 21981 8803 22015
rect 10701 21981 10735 22015
rect 12357 21981 12391 22015
rect 12633 21981 12667 22015
rect 14289 21981 14323 22015
rect 14381 21981 14415 22015
rect 15209 21981 15243 22015
rect 10149 21913 10183 21947
rect 10968 21913 11002 21947
rect 8401 21845 8435 21879
rect 8677 21845 8711 21879
rect 12081 21845 12115 21879
rect 12173 21845 12207 21879
rect 13277 21845 13311 21879
rect 14197 21845 14231 21879
rect 14473 21845 14507 21879
rect 15301 21845 15335 21879
rect 10333 21641 10367 21675
rect 6817 21505 6851 21539
rect 11161 21505 11195 21539
rect 11529 21505 11563 21539
rect 12541 21505 12575 21539
rect 12797 21505 12831 21539
rect 14381 21505 14415 21539
rect 15485 21505 15519 21539
rect 6561 21437 6595 21471
rect 8033 21437 8067 21471
rect 9413 21437 9447 21471
rect 9781 21437 9815 21471
rect 10425 21437 10459 21471
rect 11805 21437 11839 21471
rect 14565 21437 14599 21471
rect 15669 21437 15703 21471
rect 17233 21437 17267 21471
rect 18153 21437 18187 21471
rect 7941 21301 7975 21335
rect 8677 21301 8711 21335
rect 8769 21301 8803 21335
rect 11069 21301 11103 21335
rect 11253 21301 11287 21335
rect 11621 21301 11655 21335
rect 12449 21301 12483 21335
rect 13921 21301 13955 21335
rect 14289 21301 14323 21335
rect 15209 21301 15243 21335
rect 15393 21301 15427 21335
rect 16313 21301 16347 21335
rect 16681 21301 16715 21335
rect 18797 21301 18831 21335
rect 10977 21097 11011 21131
rect 15485 21097 15519 21131
rect 16957 21029 16991 21063
rect 6837 20961 6871 20995
rect 11069 20961 11103 20995
rect 14105 20961 14139 20995
rect 15577 20961 15611 20995
rect 17601 20961 17635 20995
rect 4261 20893 4295 20927
rect 4353 20893 4387 20927
rect 4537 20893 4571 20927
rect 6101 20893 6135 20927
rect 7093 20893 7127 20927
rect 8493 20893 8527 20927
rect 8585 20893 8619 20927
rect 9137 20893 9171 20927
rect 9321 20893 9355 20927
rect 9413 20893 9447 20927
rect 9597 20893 9631 20927
rect 12541 20893 12575 20927
rect 12797 20893 12831 20927
rect 14361 20893 14395 20927
rect 15844 20893 15878 20927
rect 17969 20893 18003 20927
rect 18337 20893 18371 20927
rect 19257 20893 19291 20927
rect 4804 20825 4838 20859
rect 8677 20825 8711 20859
rect 9864 20825 9898 20859
rect 11336 20825 11370 20859
rect 18889 20825 18923 20859
rect 5917 20757 5951 20791
rect 6745 20757 6779 20791
rect 8217 20757 8251 20791
rect 8401 20757 8435 20791
rect 9045 20757 9079 20791
rect 12449 20757 12483 20791
rect 13921 20757 13955 20791
rect 17049 20757 17083 20791
rect 18061 20757 18095 20791
rect 19349 20757 19383 20791
rect 9873 20553 9907 20587
rect 11345 20553 11379 20587
rect 15853 20553 15887 20587
rect 6837 20485 6871 20519
rect 8760 20485 8794 20519
rect 11796 20485 11830 20519
rect 17684 20485 17718 20519
rect 19134 20485 19168 20519
rect 4813 20417 4847 20451
rect 5080 20417 5114 20451
rect 6469 20417 6503 20451
rect 6745 20417 6779 20451
rect 8134 20417 8168 20451
rect 8493 20417 8527 20451
rect 10221 20417 10255 20451
rect 13001 20417 13035 20451
rect 13257 20417 13291 20451
rect 14473 20417 14507 20451
rect 14740 20417 14774 20451
rect 18889 20417 18923 20451
rect 8401 20349 8435 20383
rect 9965 20349 9999 20383
rect 11529 20349 11563 20383
rect 16037 20349 16071 20383
rect 17233 20349 17267 20383
rect 17417 20349 17451 20383
rect 12909 20281 12943 20315
rect 14381 20281 14415 20315
rect 16405 20281 16439 20315
rect 6193 20213 6227 20247
rect 6561 20213 6595 20247
rect 7021 20213 7055 20247
rect 16497 20213 16531 20247
rect 16681 20213 16715 20247
rect 18797 20213 18831 20247
rect 20269 20213 20303 20247
rect 5365 20009 5399 20043
rect 7021 20009 7055 20043
rect 12449 20009 12483 20043
rect 15761 20009 15795 20043
rect 9413 19941 9447 19975
rect 9597 19941 9631 19975
rect 12541 19941 12575 19975
rect 14473 19941 14507 19975
rect 4721 19873 4755 19907
rect 6745 19873 6779 19907
rect 8401 19873 8435 19907
rect 10977 19873 11011 19907
rect 8493 19805 8527 19839
rect 9045 19805 9079 19839
rect 9505 19805 9539 19839
rect 11069 19805 11103 19839
rect 13654 19805 13688 19839
rect 13921 19805 13955 19839
rect 14289 19805 14323 19839
rect 14565 19805 14599 19839
rect 15209 19805 15243 19839
rect 18521 19805 18555 19839
rect 18613 19805 18647 19839
rect 18889 19805 18923 19839
rect 19257 19805 19291 19839
rect 19524 19805 19558 19839
rect 6478 19737 6512 19771
rect 8134 19737 8168 19771
rect 9137 19737 9171 19771
rect 10732 19737 10766 19771
rect 11336 19737 11370 19771
rect 17049 19737 17083 19771
rect 18254 19737 18288 19771
rect 5273 19669 5307 19703
rect 8585 19669 8619 19703
rect 17141 19669 17175 19703
rect 18705 19669 18739 19703
rect 18981 19669 19015 19703
rect 20637 19669 20671 19703
rect 8033 19465 8067 19499
rect 16497 19465 16531 19499
rect 19809 19465 19843 19499
rect 12081 19397 12115 19431
rect 14473 19397 14507 19431
rect 14832 19397 14866 19431
rect 4721 19329 4755 19363
rect 4813 19329 4847 19363
rect 5080 19329 5114 19363
rect 6377 19329 6411 19363
rect 6469 19329 6503 19363
rect 6653 19329 6687 19363
rect 6920 19329 6954 19363
rect 8125 19329 8159 19363
rect 8392 19329 8426 19363
rect 9597 19329 9631 19363
rect 9864 19329 9898 19363
rect 11345 19329 11379 19363
rect 11621 19329 11655 19363
rect 11713 19329 11747 19363
rect 13829 19329 13863 19363
rect 17989 19329 18023 19363
rect 18337 19329 18371 19363
rect 18593 19329 18627 19363
rect 20545 19329 20579 19363
rect 23029 19329 23063 19363
rect 23305 19329 23339 19363
rect 14013 19261 14047 19295
rect 14565 19261 14599 19295
rect 16037 19261 16071 19295
rect 18245 19261 18279 19295
rect 20453 19261 20487 19295
rect 10977 19193 11011 19227
rect 14197 19193 14231 19227
rect 15945 19193 15979 19227
rect 16405 19193 16439 19227
rect 20637 19193 20671 19227
rect 4537 19125 4571 19159
rect 6193 19125 6227 19159
rect 9505 19125 9539 19159
rect 11161 19125 11195 19159
rect 16865 19125 16899 19159
rect 19717 19125 19751 19159
rect 5273 18921 5307 18955
rect 6745 18921 6779 18955
rect 8677 18921 8711 18955
rect 14197 18921 14231 18955
rect 18797 18921 18831 18955
rect 20637 18921 20671 18955
rect 8217 18853 8251 18887
rect 15945 18853 15979 18887
rect 16497 18853 16531 18887
rect 6837 18785 6871 18819
rect 11805 18785 11839 18819
rect 17877 18785 17911 18819
rect 19257 18785 19291 18819
rect 3893 18717 3927 18751
rect 4160 18717 4194 18751
rect 5365 18717 5399 18751
rect 5632 18717 5666 18751
rect 7093 18717 7127 18751
rect 8585 18717 8619 18751
rect 10517 18717 10551 18751
rect 10977 18717 11011 18751
rect 11161 18717 11195 18751
rect 13369 18717 13403 18751
rect 14105 18717 14139 18751
rect 14381 18717 14415 18751
rect 18521 18717 18555 18751
rect 18889 18717 18923 18751
rect 20729 18717 20763 18751
rect 21281 18717 21315 18751
rect 23029 18717 23063 18751
rect 8953 18649 8987 18683
rect 12072 18649 12106 18683
rect 14657 18649 14691 18683
rect 17632 18649 17666 18683
rect 19524 18649 19558 18683
rect 23305 18649 23339 18683
rect 10885 18581 10919 18615
rect 11713 18581 11747 18615
rect 13185 18581 13219 18615
rect 13921 18581 13955 18615
rect 14565 18581 14599 18615
rect 17969 18581 18003 18615
rect 4077 18377 4111 18411
rect 4353 18377 4387 18411
rect 9873 18377 9907 18411
rect 11529 18377 11563 18411
rect 15301 18377 15335 18411
rect 18061 18377 18095 18411
rect 18153 18377 18187 18411
rect 21005 18377 21039 18411
rect 6898 18309 6932 18343
rect 11345 18309 11379 18343
rect 13921 18309 13955 18343
rect 19266 18309 19300 18343
rect 19870 18309 19904 18343
rect 4169 18241 4203 18275
rect 4445 18241 4479 18275
rect 4537 18241 4571 18275
rect 5937 18241 5971 18275
rect 6193 18241 6227 18275
rect 6561 18241 6595 18275
rect 9238 18241 9272 18275
rect 12173 18241 12207 18275
rect 14013 18241 14047 18275
rect 16681 18241 16715 18275
rect 16948 18241 16982 18275
rect 6653 18173 6687 18207
rect 9505 18173 9539 18207
rect 11989 18173 12023 18207
rect 16405 18173 16439 18207
rect 19533 18173 19567 18207
rect 19625 18173 19659 18207
rect 4721 18105 4755 18139
rect 8125 18105 8159 18139
rect 11621 18105 11655 18139
rect 4813 18037 4847 18071
rect 6377 18037 6411 18071
rect 8033 18037 8067 18071
rect 15853 18037 15887 18071
rect 9137 17833 9171 17867
rect 11345 17833 11379 17867
rect 13461 17833 13495 17867
rect 14565 17833 14599 17867
rect 16129 17833 16163 17867
rect 18705 17833 18739 17867
rect 11621 17765 11655 17799
rect 14473 17765 14507 17799
rect 7021 17697 7055 17731
rect 9965 17697 9999 17731
rect 11529 17697 11563 17731
rect 12081 17697 12115 17731
rect 18429 17697 18463 17731
rect 4077 17629 4111 17663
rect 4721 17629 4755 17663
rect 6929 17629 6963 17663
rect 8953 17629 8987 17663
rect 9321 17629 9355 17663
rect 11989 17629 12023 17663
rect 13737 17629 13771 17663
rect 14105 17629 14139 17663
rect 14749 17629 14783 17663
rect 18245 17629 18279 17663
rect 18521 17629 18555 17663
rect 18797 17629 18831 17663
rect 18889 17629 18923 17663
rect 19349 17629 19383 17663
rect 4813 17561 4847 17595
rect 6561 17561 6595 17595
rect 8769 17561 8803 17595
rect 10210 17561 10244 17595
rect 12326 17561 12360 17595
rect 14994 17561 15028 17595
rect 16221 17561 16255 17595
rect 6837 17493 6871 17527
rect 9873 17493 9907 17527
rect 13645 17493 13679 17527
rect 17509 17493 17543 17527
rect 18153 17493 18187 17527
rect 18981 17493 19015 17527
rect 19441 17493 19475 17527
rect 4721 17289 4755 17323
rect 6745 17289 6779 17323
rect 10885 17289 10919 17323
rect 11529 17289 11563 17323
rect 13277 17289 13311 17323
rect 14749 17289 14783 17323
rect 16405 17289 16439 17323
rect 17969 17289 18003 17323
rect 7481 17221 7515 17255
rect 9229 17221 9263 17255
rect 12164 17221 12198 17255
rect 1869 17153 1903 17187
rect 3433 17153 3467 17187
rect 3709 17153 3743 17187
rect 3985 17153 4019 17187
rect 4813 17153 4847 17187
rect 5080 17153 5114 17187
rect 6469 17153 6503 17187
rect 9321 17153 9355 17187
rect 9597 17153 9631 17187
rect 11713 17153 11747 17187
rect 13369 17153 13403 17187
rect 13636 17153 13670 17187
rect 15025 17153 15059 17187
rect 15292 17153 15326 17187
rect 16681 17153 16715 17187
rect 19634 17153 19668 17187
rect 19993 17153 20027 17187
rect 20260 17153 20294 17187
rect 23029 17153 23063 17187
rect 1593 17085 1627 17119
rect 4169 17085 4203 17119
rect 7297 17085 7331 17119
rect 11897 17085 11931 17119
rect 19901 17085 19935 17119
rect 23305 17085 23339 17119
rect 3617 17017 3651 17051
rect 6561 17017 6595 17051
rect 21373 17017 21407 17051
rect 3249 16949 3283 16983
rect 3893 16949 3927 16983
rect 6193 16949 6227 16983
rect 9413 16949 9447 16983
rect 18521 16949 18555 16983
rect 6745 16745 6779 16779
rect 11621 16745 11655 16779
rect 21189 16745 21223 16779
rect 8401 16677 8435 16711
rect 9045 16677 9079 16711
rect 12357 16677 12391 16711
rect 18705 16677 18739 16711
rect 3065 16609 3099 16643
rect 6377 16609 6411 16643
rect 12265 16609 12299 16643
rect 13737 16609 13771 16643
rect 17693 16609 17727 16643
rect 21097 16609 21131 16643
rect 22477 16609 22511 16643
rect 2145 16541 2179 16575
rect 2697 16541 2731 16575
rect 3985 16541 4019 16575
rect 4353 16541 4387 16575
rect 6121 16541 6155 16575
rect 11345 16541 11379 16575
rect 13470 16541 13504 16575
rect 15853 16541 15887 16575
rect 18429 16541 18463 16575
rect 19257 16541 19291 16575
rect 21741 16541 21775 16575
rect 22845 16541 22879 16575
rect 23029 16541 23063 16575
rect 2789 16473 2823 16507
rect 4905 16473 4939 16507
rect 8217 16473 8251 16507
rect 8769 16473 8803 16507
rect 9413 16473 9447 16507
rect 14105 16473 14139 16507
rect 15945 16473 15979 16507
rect 18981 16473 19015 16507
rect 20830 16473 20864 16507
rect 23305 16473 23339 16507
rect 2053 16405 2087 16439
rect 3617 16405 3651 16439
rect 4077 16405 4111 16439
rect 4997 16405 5031 16439
rect 8309 16405 8343 16439
rect 8953 16405 8987 16439
rect 9873 16405 9907 16439
rect 17785 16405 17819 16439
rect 18521 16405 18555 16439
rect 19349 16405 19383 16439
rect 19717 16405 19751 16439
rect 21925 16405 21959 16439
rect 22753 16405 22787 16439
rect 3341 16201 3375 16235
rect 6193 16201 6227 16235
rect 6561 16201 6595 16235
rect 11529 16201 11563 16235
rect 12081 16201 12115 16235
rect 14381 16201 14415 16235
rect 18429 16201 18463 16235
rect 20637 16201 20671 16235
rect 5058 16133 5092 16167
rect 10609 16133 10643 16167
rect 11989 16133 12023 16167
rect 13194 16133 13228 16167
rect 16957 16133 16991 16167
rect 18797 16133 18831 16167
rect 1869 16065 1903 16099
rect 2053 16065 2087 16099
rect 2329 16065 2363 16099
rect 2697 16065 2731 16099
rect 4454 16065 4488 16099
rect 4813 16065 4847 16099
rect 6653 16065 6687 16099
rect 7858 16065 7892 16099
rect 8125 16065 8159 16099
rect 8217 16065 8251 16099
rect 13461 16065 13495 16099
rect 14473 16065 14507 16099
rect 15016 16065 15050 16099
rect 16221 16065 16255 16099
rect 16681 16065 16715 16099
rect 21557 16065 21591 16099
rect 22017 16065 22051 16099
rect 1593 15997 1627 16031
rect 2145 15997 2179 16031
rect 4721 15997 4755 16031
rect 11345 15997 11379 16031
rect 14105 15997 14139 16031
rect 14749 15997 14783 16031
rect 21189 15997 21223 16031
rect 22109 15997 22143 16031
rect 23397 15997 23431 16031
rect 9505 15929 9539 15963
rect 10333 15929 10367 15963
rect 10701 15929 10735 15963
rect 11713 15929 11747 15963
rect 20085 15929 20119 15963
rect 21925 15929 21959 15963
rect 2513 15861 2547 15895
rect 3249 15861 3283 15895
rect 6745 15861 6779 15895
rect 10149 15861 10183 15895
rect 13553 15861 13587 15895
rect 16129 15861 16163 15895
rect 16313 15861 16347 15895
rect 16773 15861 16807 15895
rect 21465 15861 21499 15895
rect 22753 15861 22787 15895
rect 22845 15861 22879 15895
rect 1685 15657 1719 15691
rect 3617 15657 3651 15691
rect 3985 15657 4019 15691
rect 7297 15657 7331 15691
rect 7389 15657 7423 15691
rect 11989 15657 12023 15691
rect 13461 15657 13495 15691
rect 14381 15657 14415 15691
rect 5825 15589 5859 15623
rect 20545 15589 20579 15623
rect 4445 15521 4479 15555
rect 8769 15521 8803 15555
rect 10609 15521 10643 15555
rect 17693 15521 17727 15555
rect 22477 15521 22511 15555
rect 23397 15521 23431 15555
rect 1593 15453 1627 15487
rect 2053 15453 2087 15487
rect 2329 15453 2363 15487
rect 2605 15453 2639 15487
rect 2697 15453 2731 15487
rect 3065 15453 3099 15487
rect 4077 15453 4111 15487
rect 4169 15453 4203 15487
rect 5917 15453 5951 15487
rect 10425 15453 10459 15487
rect 10876 15453 10910 15487
rect 12081 15453 12115 15487
rect 13921 15453 13955 15487
rect 14289 15453 14323 15487
rect 15761 15453 15795 15487
rect 17601 15453 17635 15487
rect 19257 15453 19291 15487
rect 22221 15453 22255 15487
rect 23121 15453 23155 15487
rect 23305 15453 23339 15487
rect 2513 15385 2547 15419
rect 4261 15385 4295 15419
rect 4712 15385 4746 15419
rect 6162 15385 6196 15419
rect 8502 15385 8536 15419
rect 10158 15385 10192 15419
rect 12348 15385 12382 15419
rect 14197 15385 14231 15419
rect 15516 15385 15550 15419
rect 15853 15385 15887 15419
rect 17960 15385 17994 15419
rect 1961 15317 1995 15351
rect 2145 15317 2179 15351
rect 2789 15317 2823 15351
rect 9045 15317 9079 15351
rect 13829 15317 13863 15351
rect 19073 15317 19107 15351
rect 21097 15317 21131 15351
rect 22569 15317 22603 15351
rect 6193 15113 6227 15147
rect 7757 15113 7791 15147
rect 8309 15113 8343 15147
rect 9781 15113 9815 15147
rect 12357 15113 12391 15147
rect 14381 15113 14415 15147
rect 21833 15113 21867 15147
rect 2136 15045 2170 15079
rect 13492 15045 13526 15079
rect 15669 15045 15703 15079
rect 19870 15045 19904 15079
rect 1593 14977 1627 15011
rect 3341 14977 3375 15011
rect 3597 14977 3631 15011
rect 4813 14977 4847 15011
rect 5069 14977 5103 15011
rect 6377 14977 6411 15011
rect 6633 14977 6667 15011
rect 9597 14977 9631 15011
rect 9689 14977 9723 15011
rect 9965 14977 9999 15011
rect 10232 14977 10266 15011
rect 12265 14977 12299 15011
rect 13737 14977 13771 15011
rect 16681 14977 16715 15011
rect 16948 14977 16982 15011
rect 18153 14977 18187 15011
rect 18409 14977 18443 15011
rect 19625 14977 19659 15011
rect 21097 14977 21131 15011
rect 21557 14977 21591 15011
rect 22957 14977 22991 15011
rect 23213 14977 23247 15011
rect 23305 14977 23339 15011
rect 1869 14909 1903 14943
rect 16313 14909 16347 14943
rect 3249 14841 3283 14875
rect 4721 14841 4755 14875
rect 21005 14841 21039 14875
rect 1685 14773 1719 14807
rect 11345 14773 11379 14807
rect 11621 14773 11655 14807
rect 15761 14773 15795 14807
rect 18061 14773 18095 14807
rect 19533 14773 19567 14807
rect 21189 14773 21223 14807
rect 21465 14773 21499 14807
rect 23397 14773 23431 14807
rect 17049 14569 17083 14603
rect 3617 14501 3651 14535
rect 5273 14501 5307 14535
rect 5365 14501 5399 14535
rect 18889 14501 18923 14535
rect 20637 14501 20671 14535
rect 2329 14433 2363 14467
rect 3893 14433 3927 14467
rect 6745 14433 6779 14467
rect 9597 14433 9631 14467
rect 13093 14433 13127 14467
rect 14105 14433 14139 14467
rect 15577 14433 15611 14467
rect 18429 14433 18463 14467
rect 18521 14433 18555 14467
rect 2053 14365 2087 14399
rect 3065 14365 3099 14399
rect 6478 14365 6512 14399
rect 9689 14365 9723 14399
rect 13185 14365 13219 14399
rect 13369 14365 13403 14399
rect 13921 14365 13955 14399
rect 14361 14365 14395 14399
rect 15833 14365 15867 14399
rect 18162 14365 18196 14399
rect 19257 14365 19291 14399
rect 22109 14365 22143 14399
rect 22753 14365 22787 14399
rect 23029 14365 23063 14399
rect 1501 14297 1535 14331
rect 2881 14297 2915 14331
rect 4160 14297 4194 14331
rect 8585 14297 8619 14331
rect 9956 14297 9990 14331
rect 12909 14297 12943 14331
rect 19524 14297 19558 14331
rect 21864 14297 21898 14331
rect 23305 14297 23339 14331
rect 7113 14229 7147 14263
rect 8953 14229 8987 14263
rect 11069 14229 11103 14263
rect 11437 14229 11471 14263
rect 15485 14229 15519 14263
rect 16957 14229 16991 14263
rect 18981 14229 19015 14263
rect 20729 14229 20763 14263
rect 22201 14229 22235 14263
rect 1777 14025 1811 14059
rect 13461 14025 13495 14059
rect 15393 14025 15427 14059
rect 16497 14025 16531 14059
rect 16865 14025 16899 14059
rect 16957 14025 16991 14059
rect 17693 14025 17727 14059
rect 20637 14025 20671 14059
rect 23397 14025 23431 14059
rect 7604 13957 7638 13991
rect 11529 13957 11563 13991
rect 13553 13957 13587 13991
rect 18806 13957 18840 13991
rect 1593 13889 1627 13923
rect 1869 13889 1903 13923
rect 2136 13889 2170 13923
rect 3341 13889 3375 13923
rect 3597 13889 3631 13923
rect 5080 13889 5114 13923
rect 7849 13889 7883 13923
rect 7941 13889 7975 13923
rect 11078 13889 11112 13923
rect 12081 13889 12115 13923
rect 12337 13889 12371 13923
rect 15577 13889 15611 13923
rect 15945 13889 15979 13923
rect 16681 13889 16715 13923
rect 17509 13889 17543 13923
rect 19073 13889 19107 13923
rect 20289 13889 20323 13923
rect 20545 13889 20579 13923
rect 21557 13889 21591 13923
rect 21833 13889 21867 13923
rect 22100 13889 22134 13923
rect 23305 13879 23339 13913
rect 4813 13821 4847 13855
rect 9505 13821 9539 13855
rect 11345 13821 11379 13855
rect 11989 13821 12023 13855
rect 21281 13821 21315 13855
rect 3249 13753 3283 13787
rect 4721 13753 4755 13787
rect 6193 13753 6227 13787
rect 6469 13753 6503 13787
rect 9965 13753 9999 13787
rect 11805 13753 11839 13787
rect 19165 13753 19199 13787
rect 23213 13753 23247 13787
rect 14841 13685 14875 13719
rect 21373 13685 21407 13719
rect 10793 13481 10827 13515
rect 13553 13481 13587 13515
rect 16773 13481 16807 13515
rect 18705 13481 18739 13515
rect 22109 13481 22143 13515
rect 3893 13413 3927 13447
rect 7297 13413 7331 13447
rect 13829 13413 13863 13447
rect 14289 13413 14323 13447
rect 1501 13345 1535 13379
rect 4077 13345 4111 13379
rect 13185 13345 13219 13379
rect 23397 13345 23431 13379
rect 2053 13277 2087 13311
rect 3617 13277 3651 13311
rect 3801 13277 3835 13311
rect 5549 13277 5583 13311
rect 10701 13277 10735 13311
rect 11345 13277 11379 13311
rect 11621 13277 11655 13311
rect 13461 13277 13495 13311
rect 13921 13277 13955 13311
rect 14105 13277 14139 13311
rect 14381 13277 14415 13311
rect 14749 13277 14783 13311
rect 17325 13277 17359 13311
rect 18981 13277 19015 13311
rect 20637 13277 20671 13311
rect 20729 13277 20763 13311
rect 22201 13277 22235 13311
rect 22845 13277 22879 13311
rect 3350 13209 3384 13243
rect 4344 13209 4378 13243
rect 5816 13209 5850 13243
rect 8769 13209 8803 13243
rect 15485 13209 15519 13243
rect 17592 13209 17626 13243
rect 20392 13209 20426 13243
rect 20996 13209 21030 13243
rect 22477 13209 22511 13243
rect 2237 13141 2271 13175
rect 5457 13141 5491 13175
rect 6929 13141 6963 13175
rect 9413 13141 9447 13175
rect 14565 13141 14599 13175
rect 15393 13141 15427 13175
rect 18889 13141 18923 13175
rect 19257 13141 19291 13175
rect 1685 12937 1719 12971
rect 6469 12937 6503 12971
rect 12817 12937 12851 12971
rect 13829 12937 13863 12971
rect 18337 12937 18371 12971
rect 19809 12937 19843 12971
rect 6745 12869 6779 12903
rect 10885 12869 10919 12903
rect 22100 12869 22134 12903
rect 1777 12801 1811 12835
rect 2993 12801 3027 12835
rect 3249 12801 3283 12835
rect 3341 12801 3375 12835
rect 3597 12801 3631 12835
rect 5069 12801 5103 12835
rect 6377 12801 6411 12835
rect 6837 12801 6871 12835
rect 7021 12801 7055 12835
rect 7665 12801 7699 12835
rect 7921 12801 7955 12835
rect 11345 12801 11379 12835
rect 11529 12801 11563 12835
rect 13553 12801 13587 12835
rect 13645 12801 13679 12835
rect 13921 12801 13955 12835
rect 15597 12801 15631 12835
rect 15853 12801 15887 12835
rect 15945 12801 15979 12835
rect 16865 12801 16899 12835
rect 17132 12801 17166 12835
rect 19461 12801 19495 12835
rect 20922 12801 20956 12835
rect 21465 12801 21499 12835
rect 23305 12801 23339 12835
rect 4813 12733 4847 12767
rect 19717 12733 19751 12767
rect 21189 12733 21223 12767
rect 21833 12733 21867 12767
rect 23397 12733 23431 12767
rect 14289 12665 14323 12699
rect 14473 12665 14507 12699
rect 16221 12665 16255 12699
rect 18245 12665 18279 12699
rect 1869 12597 1903 12631
rect 4721 12597 4755 12631
rect 6193 12597 6227 12631
rect 7573 12597 7607 12631
rect 9045 12597 9079 12631
rect 9597 12597 9631 12631
rect 11161 12597 11195 12631
rect 13461 12597 13495 12631
rect 14381 12597 14415 12631
rect 16405 12597 16439 12631
rect 21373 12597 21407 12631
rect 23213 12597 23247 12631
rect 3617 12393 3651 12427
rect 13737 12393 13771 12427
rect 22661 12393 22695 12427
rect 11621 12325 11655 12359
rect 12081 12325 12115 12359
rect 18889 12325 18923 12359
rect 2237 12257 2271 12291
rect 4353 12257 4387 12291
rect 8769 12257 8803 12291
rect 13461 12257 13495 12291
rect 1501 12189 1535 12223
rect 2053 12189 2087 12223
rect 7297 12189 7331 12223
rect 8513 12189 8547 12223
rect 8953 12189 8987 12223
rect 10793 12189 10827 12223
rect 11345 12189 11379 12223
rect 13205 12189 13239 12223
rect 13553 12189 13587 12223
rect 15229 12189 15263 12223
rect 15485 12189 15519 12223
rect 15669 12189 15703 12223
rect 15761 12189 15795 12223
rect 16037 12189 16071 12223
rect 17969 12189 18003 12223
rect 18521 12189 18555 12223
rect 18797 12189 18831 12223
rect 19073 12189 19107 12223
rect 19257 12189 19291 12223
rect 2504 12121 2538 12155
rect 4598 12121 4632 12155
rect 7052 12121 7086 12155
rect 11989 12121 12023 12155
rect 21189 12121 21223 12155
rect 5733 12053 5767 12087
rect 5917 12053 5951 12087
rect 7389 12053 7423 12087
rect 10241 12053 10275 12087
rect 11529 12053 11563 12087
rect 14105 12053 14139 12087
rect 17325 12053 17359 12087
rect 18613 12053 18647 12087
rect 20545 12053 20579 12087
rect 11161 11849 11195 11883
rect 21557 11849 21591 11883
rect 23397 11849 23431 11883
rect 2114 11781 2148 11815
rect 7849 11781 7883 11815
rect 9934 11781 9968 11815
rect 13093 11781 13127 11815
rect 14841 11781 14875 11815
rect 18429 11781 18463 11815
rect 22100 11781 22134 11815
rect 1593 11713 1627 11747
rect 3597 11713 3631 11747
rect 5937 11713 5971 11747
rect 6193 11713 6227 11747
rect 6644 11713 6678 11747
rect 9689 11713 9723 11747
rect 11345 11713 11379 11747
rect 11621 11713 11655 11747
rect 11877 11713 11911 11747
rect 15200 11713 15234 11747
rect 18521 11713 18555 11747
rect 18777 11713 18811 11747
rect 21117 11713 21151 11747
rect 21649 11713 21683 11747
rect 23305 11713 23339 11747
rect 1869 11645 1903 11679
rect 3341 11645 3375 11679
rect 6377 11645 6411 11679
rect 14933 11645 14967 11679
rect 21373 11645 21407 11679
rect 21833 11645 21867 11679
rect 1777 11577 1811 11611
rect 4813 11577 4847 11611
rect 11069 11577 11103 11611
rect 16313 11577 16347 11611
rect 23213 11577 23247 11611
rect 3249 11509 3283 11543
rect 4721 11509 4755 11543
rect 7757 11509 7791 11543
rect 9137 11509 9171 11543
rect 13001 11509 13035 11543
rect 16957 11509 16991 11543
rect 19901 11509 19935 11543
rect 19993 11509 20027 11543
rect 2145 11305 2179 11339
rect 5825 11305 5859 11339
rect 8769 11305 8803 11339
rect 12173 11305 12207 11339
rect 13829 11305 13863 11339
rect 11253 11237 11287 11271
rect 15301 11237 15335 11271
rect 16773 11237 16807 11271
rect 19625 11237 19659 11271
rect 11345 11169 11379 11203
rect 11989 11169 12023 11203
rect 13553 11169 13587 11203
rect 14657 11169 14691 11203
rect 17141 11169 17175 11203
rect 19257 11169 19291 11203
rect 19717 11169 19751 11203
rect 21557 11169 21591 11203
rect 1593 11101 1627 11135
rect 2237 11101 2271 11135
rect 4445 11101 4479 11135
rect 6101 11101 6135 11135
rect 7389 11101 7423 11135
rect 7656 11101 7690 11135
rect 11437 11101 11471 11135
rect 13286 11101 13320 11135
rect 13645 11101 13679 11135
rect 16589 11101 16623 11135
rect 18889 11101 18923 11135
rect 19809 11101 19843 11135
rect 23029 11101 23063 11135
rect 23121 11101 23155 11135
rect 23213 11101 23247 11135
rect 2504 11033 2538 11067
rect 4690 11033 4724 11067
rect 6469 11033 6503 11067
rect 8953 11033 8987 11067
rect 10517 11033 10551 11067
rect 10885 11033 10919 11067
rect 14105 11033 14139 11067
rect 17325 11033 17359 11067
rect 22762 11033 22796 11067
rect 3617 10965 3651 10999
rect 16681 10965 16715 10999
rect 21649 10965 21683 10999
rect 4629 10761 4663 10795
rect 15485 10761 15519 10795
rect 16221 10761 16255 10795
rect 16773 10761 16807 10795
rect 21097 10761 21131 10795
rect 23397 10761 23431 10795
rect 8493 10693 8527 10727
rect 1501 10625 1535 10659
rect 2033 10625 2067 10659
rect 3249 10625 3283 10659
rect 3505 10625 3539 10659
rect 5069 10625 5103 10659
rect 6469 10625 6503 10659
rect 8585 10625 8619 10659
rect 11161 10625 11195 10659
rect 11621 10625 11655 10659
rect 13481 10625 13515 10659
rect 13737 10625 13771 10659
rect 14013 10625 14047 10659
rect 14372 10625 14406 10659
rect 15577 10625 15611 10659
rect 16313 10625 16347 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 18797 10625 18831 10659
rect 20013 10625 20047 10659
rect 21281 10625 21315 10659
rect 21373 10625 21407 10659
rect 22946 10625 22980 10659
rect 23213 10625 23247 10659
rect 23305 10625 23339 10659
rect 1777 10557 1811 10591
rect 4813 10557 4847 10591
rect 11069 10557 11103 10591
rect 12265 10557 12299 10591
rect 14105 10557 14139 10591
rect 20269 10557 20303 10591
rect 21005 10557 21039 10591
rect 3157 10489 3191 10523
rect 6193 10489 6227 10523
rect 6653 10489 6687 10523
rect 11345 10489 11379 10523
rect 12357 10489 12391 10523
rect 16405 10489 16439 10523
rect 21465 10489 21499 10523
rect 21833 10489 21867 10523
rect 1685 10421 1719 10455
rect 7021 10421 7055 10455
rect 10057 10421 10091 10455
rect 10425 10421 10459 10455
rect 13921 10421 13955 10455
rect 18889 10421 18923 10455
rect 20361 10421 20395 10455
rect 6009 10217 6043 10251
rect 8125 10217 8159 10251
rect 12265 10217 12299 10251
rect 13921 10217 13955 10251
rect 15669 10217 15703 10251
rect 20637 10217 20671 10251
rect 3617 10149 3651 10183
rect 9137 10149 9171 10183
rect 18797 10149 18831 10183
rect 1593 10081 1627 10115
rect 3985 10081 4019 10115
rect 8769 10081 8803 10115
rect 18521 10081 18555 10115
rect 23305 10081 23339 10115
rect 2881 10013 2915 10047
rect 3065 10013 3099 10047
rect 5733 10013 5767 10047
rect 5917 10013 5951 10047
rect 9505 10013 9539 10047
rect 11897 10013 11931 10047
rect 12081 10013 12115 10047
rect 12541 10013 12575 10047
rect 12808 10013 12842 10047
rect 15577 10013 15611 10047
rect 17049 10013 17083 10047
rect 19257 10013 19291 10047
rect 20729 10013 20763 10047
rect 22201 10013 22235 10047
rect 22477 10013 22511 10047
rect 22845 10013 22879 10047
rect 2145 9945 2179 9979
rect 6193 9945 6227 9979
rect 7941 9945 7975 9979
rect 9413 9945 9447 9979
rect 15310 9945 15344 9979
rect 16804 9945 16838 9979
rect 18254 9945 18288 9979
rect 19073 9945 19107 9979
rect 19502 9945 19536 9979
rect 20996 9945 21030 9979
rect 2237 9877 2271 9911
rect 8953 9877 8987 9911
rect 10793 9877 10827 9911
rect 11345 9877 11379 9911
rect 14197 9877 14231 9911
rect 17141 9877 17175 9911
rect 18613 9877 18647 9911
rect 22109 9877 22143 9911
rect 2145 9605 2179 9639
rect 6377 9605 6411 9639
rect 13952 9605 13986 9639
rect 14657 9605 14691 9639
rect 16405 9605 16439 9639
rect 16681 9605 16715 9639
rect 19634 9605 19668 9639
rect 21106 9605 21140 9639
rect 2237 9537 2271 9571
rect 2697 9537 2731 9571
rect 3249 9537 3283 9571
rect 4465 9537 4499 9571
rect 4721 9537 4755 9571
rect 5069 9537 5103 9571
rect 8125 9537 8159 9571
rect 10517 9537 10551 9571
rect 10609 9537 10643 9571
rect 11805 9537 11839 9571
rect 14473 9537 14507 9571
rect 19901 9537 19935 9571
rect 21465 9537 21499 9571
rect 22089 9537 22123 9571
rect 23489 9537 23523 9571
rect 1593 9469 1627 9503
rect 4813 9469 4847 9503
rect 8217 9469 8251 9503
rect 8677 9469 8711 9503
rect 11253 9469 11287 9503
rect 12541 9469 12575 9503
rect 14197 9469 14231 9503
rect 14381 9469 14415 9503
rect 21366 9469 21400 9503
rect 21833 9469 21867 9503
rect 2421 9401 2455 9435
rect 8401 9401 8435 9435
rect 18521 9401 18555 9435
rect 19993 9401 20027 9435
rect 21557 9401 21591 9435
rect 23305 9401 23339 9435
rect 3341 9333 3375 9367
rect 6193 9333 6227 9367
rect 9229 9333 9263 9367
rect 11621 9333 11655 9367
rect 11989 9333 12023 9367
rect 12817 9333 12851 9367
rect 17969 9333 18003 9367
rect 23213 9333 23247 9367
rect 2145 9129 2179 9163
rect 9045 9129 9079 9163
rect 10609 9129 10643 9163
rect 11989 9129 12023 9163
rect 12541 9129 12575 9163
rect 17417 9129 17451 9163
rect 18429 9061 18463 9095
rect 18889 9061 18923 9095
rect 20637 9061 20671 9095
rect 17785 8993 17819 9027
rect 23121 8993 23155 9027
rect 1593 8925 1627 8959
rect 2237 8925 2271 8959
rect 3801 8925 3835 8959
rect 4077 8925 4111 8959
rect 8769 8925 8803 8959
rect 9137 8925 9171 8959
rect 9229 8925 9263 8959
rect 10701 8925 10735 8959
rect 13921 8925 13955 8959
rect 15853 8925 15887 8959
rect 19257 8925 19291 8959
rect 20729 8925 20763 8959
rect 22845 8925 22879 8959
rect 2482 8857 2516 8891
rect 4344 8857 4378 8891
rect 7021 8857 7055 8891
rect 9496 8857 9530 8891
rect 13654 8857 13688 8891
rect 14105 8857 14139 8891
rect 15945 8857 15979 8891
rect 18521 8857 18555 8891
rect 19502 8857 19536 8891
rect 20974 8857 21008 8891
rect 3617 8789 3651 8823
rect 3985 8789 4019 8823
rect 5457 8789 5491 8823
rect 18981 8789 19015 8823
rect 22109 8789 22143 8823
rect 1685 8585 1719 8619
rect 14381 8585 14415 8619
rect 16221 8585 16255 8619
rect 19257 8585 19291 8619
rect 21373 8585 21407 8619
rect 23213 8585 23247 8619
rect 3608 8517 3642 8551
rect 6377 8517 6411 8551
rect 7941 8517 7975 8551
rect 9413 8517 9447 8551
rect 11345 8517 11379 8551
rect 14197 8517 14231 8551
rect 17417 8517 17451 8551
rect 20922 8517 20956 8551
rect 23397 8517 23431 8551
rect 1777 8449 1811 8483
rect 2993 8449 3027 8483
rect 5937 8449 5971 8483
rect 8217 8449 8251 8483
rect 12449 8449 12483 8483
rect 14473 8449 14507 8483
rect 15770 8449 15804 8483
rect 16313 8449 16347 8483
rect 16773 8449 16807 8483
rect 17325 8449 17359 8483
rect 17969 8449 18003 8483
rect 21189 8449 21223 8483
rect 21281 8449 21315 8483
rect 21833 8449 21867 8483
rect 22089 8449 22123 8483
rect 23305 8449 23339 8483
rect 3249 8381 3283 8415
rect 3341 8381 3375 8415
rect 6193 8381 6227 8415
rect 11805 8381 11839 8415
rect 16037 8381 16071 8415
rect 1869 8313 1903 8347
rect 8861 8313 8895 8347
rect 9045 8313 9079 8347
rect 12357 8313 12391 8347
rect 14657 8313 14691 8347
rect 17785 8313 17819 8347
rect 17877 8313 17911 8347
rect 4721 8245 4755 8279
rect 4813 8245 4847 8279
rect 8953 8245 8987 8279
rect 10057 8245 10091 8279
rect 19809 8245 19843 8279
rect 3617 8041 3651 8075
rect 3985 8041 4019 8075
rect 8953 8041 8987 8075
rect 12265 8041 12299 8075
rect 23213 8041 23247 8075
rect 4077 7973 4111 8007
rect 10425 7973 10459 8007
rect 10701 7905 10735 7939
rect 19809 7905 19843 7939
rect 1593 7837 1627 7871
rect 2237 7837 2271 7871
rect 3801 7837 3835 7871
rect 5457 7837 5491 7871
rect 5549 7837 5583 7871
rect 5805 7837 5839 7871
rect 7389 7837 7423 7871
rect 10333 7837 10367 7871
rect 10609 7837 10643 7871
rect 12173 7837 12207 7871
rect 13921 7837 13955 7871
rect 14197 7837 14231 7871
rect 14289 7837 14323 7871
rect 15945 7837 15979 7871
rect 16037 7837 16071 7871
rect 18889 7837 18923 7871
rect 21557 7837 21591 7871
rect 23029 7837 23063 7871
rect 23305 7837 23339 7871
rect 2504 7769 2538 7803
rect 5190 7769 5224 7803
rect 7634 7769 7668 7803
rect 10066 7769 10100 7803
rect 10968 7769 11002 7803
rect 13654 7769 13688 7803
rect 15700 7769 15734 7803
rect 16304 7769 16338 7803
rect 18622 7769 18656 7803
rect 19257 7769 19291 7803
rect 21312 7769 21346 7803
rect 22762 7769 22796 7803
rect 2145 7701 2179 7735
rect 6929 7701 6963 7735
rect 8769 7701 8803 7735
rect 12081 7701 12115 7735
rect 12541 7701 12575 7735
rect 14565 7701 14599 7735
rect 17417 7701 17451 7735
rect 17509 7701 17543 7735
rect 20177 7701 20211 7735
rect 21649 7701 21683 7735
rect 2421 7497 2455 7531
rect 9873 7497 9907 7531
rect 12081 7497 12115 7531
rect 13553 7497 13587 7531
rect 14749 7497 14783 7531
rect 16313 7497 16347 7531
rect 21465 7497 21499 7531
rect 2053 7429 2087 7463
rect 3249 7429 3283 7463
rect 3586 7429 3620 7463
rect 8738 7429 8772 7463
rect 14473 7429 14507 7463
rect 1777 7361 1811 7395
rect 1961 7361 1995 7395
rect 2513 7361 2547 7395
rect 5926 7361 5960 7395
rect 7021 7361 7055 7395
rect 7288 7361 7322 7395
rect 11089 7361 11123 7395
rect 11345 7361 11379 7395
rect 12429 7361 12463 7395
rect 13645 7361 13679 7395
rect 14381 7361 14415 7395
rect 15862 7361 15896 7395
rect 16129 7361 16163 7395
rect 16221 7361 16255 7395
rect 17805 7361 17839 7395
rect 19266 7361 19300 7395
rect 19533 7361 19567 7395
rect 19881 7361 19915 7395
rect 21281 7361 21315 7395
rect 21557 7361 21591 7395
rect 22957 7361 22991 7395
rect 23297 7351 23331 7385
rect 2697 7293 2731 7327
rect 3341 7293 3375 7327
rect 6193 7293 6227 7327
rect 6929 7293 6963 7327
rect 8493 7293 8527 7327
rect 11621 7293 11655 7327
rect 12173 7293 12207 7327
rect 14289 7293 14323 7327
rect 18061 7293 18095 7327
rect 19625 7293 19659 7327
rect 21189 7293 21223 7327
rect 23213 7293 23247 7327
rect 1685 7225 1719 7259
rect 4813 7225 4847 7259
rect 6653 7225 6687 7259
rect 11897 7225 11931 7259
rect 18153 7225 18187 7259
rect 21005 7225 21039 7259
rect 23397 7225 23431 7259
rect 4721 7157 4755 7191
rect 6469 7157 6503 7191
rect 8401 7157 8435 7191
rect 9965 7157 9999 7191
rect 16681 7157 16715 7191
rect 21833 7157 21867 7191
rect 1593 6953 1627 6987
rect 2053 6953 2087 6987
rect 3893 6953 3927 6987
rect 15485 6953 15519 6987
rect 18797 6953 18831 6987
rect 9045 6885 9079 6919
rect 9229 6885 9263 6919
rect 1777 6817 1811 6851
rect 2789 6817 2823 6851
rect 2973 6817 3007 6851
rect 4169 6817 4203 6851
rect 9597 6817 9631 6851
rect 23121 6817 23155 6851
rect 1409 6749 1443 6783
rect 1869 6749 1903 6783
rect 1961 6749 1995 6783
rect 2605 6749 2639 6783
rect 2881 6749 2915 6783
rect 3801 6749 3835 6783
rect 4077 6749 4111 6783
rect 4353 6749 4387 6783
rect 7297 6749 7331 6783
rect 11069 6749 11103 6783
rect 14105 6749 14139 6783
rect 14372 6749 14406 6783
rect 16957 6749 16991 6783
rect 17233 6749 17267 6783
rect 18889 6749 18923 6783
rect 19257 6749 19291 6783
rect 20729 6749 20763 6783
rect 22845 6749 22879 6783
rect 4598 6681 4632 6715
rect 7564 6681 7598 6715
rect 9505 6681 9539 6715
rect 9864 6681 9898 6715
rect 11336 6681 11370 6715
rect 16712 6681 16746 6715
rect 17500 6681 17534 6715
rect 19524 6681 19558 6715
rect 20996 6681 21030 6715
rect 2513 6613 2547 6647
rect 3617 6613 3651 6647
rect 5733 6613 5767 6647
rect 8677 6613 8711 6647
rect 10977 6613 11011 6647
rect 12449 6613 12483 6647
rect 15577 6613 15611 6647
rect 18613 6613 18647 6647
rect 20637 6613 20671 6647
rect 22109 6613 22143 6647
rect 1685 6409 1719 6443
rect 4721 6409 4755 6443
rect 6561 6409 6595 6443
rect 6837 6409 6871 6443
rect 9873 6409 9907 6443
rect 11529 6409 11563 6443
rect 12541 6409 12575 6443
rect 16405 6409 16439 6443
rect 16773 6409 16807 6443
rect 18521 6409 18555 6443
rect 21281 6409 21315 6443
rect 23397 6409 23431 6443
rect 14350 6341 14384 6375
rect 20116 6341 20150 6375
rect 1777 6273 1811 6307
rect 2136 6273 2170 6307
rect 3341 6273 3375 6307
rect 3608 6273 3642 6307
rect 5069 6273 5103 6307
rect 6653 6273 6687 6307
rect 6929 6273 6963 6307
rect 7277 6273 7311 6307
rect 8493 6273 8527 6307
rect 8760 6273 8794 6307
rect 9965 6273 9999 6307
rect 10232 6273 10266 6307
rect 12081 6273 12115 6307
rect 13654 6273 13688 6307
rect 13921 6273 13955 6307
rect 16129 6273 16163 6307
rect 16497 6273 16531 6307
rect 16865 6273 16899 6307
rect 18162 6273 18196 6307
rect 18705 6273 18739 6307
rect 20453 6273 20487 6307
rect 21097 6273 21131 6307
rect 21373 6273 21407 6307
rect 21649 6273 21683 6307
rect 22957 6273 22991 6307
rect 23305 6273 23339 6307
rect 1869 6205 1903 6239
rect 4813 6205 4847 6239
rect 7021 6205 7055 6239
rect 14105 6205 14139 6239
rect 18429 6205 18463 6239
rect 20361 6205 20395 6239
rect 23213 6205 23247 6239
rect 21557 6137 21591 6171
rect 3249 6069 3283 6103
rect 6193 6069 6227 6103
rect 8401 6069 8435 6103
rect 11345 6069 11379 6103
rect 15485 6069 15519 6103
rect 15577 6069 15611 6103
rect 17049 6069 17083 6103
rect 18981 6069 19015 6103
rect 21833 6069 21867 6103
rect 2329 5865 2363 5899
rect 2881 5865 2915 5899
rect 3893 5865 3927 5899
rect 4169 5865 4203 5899
rect 9045 5865 9079 5899
rect 14657 5865 14691 5899
rect 18981 5865 19015 5899
rect 19349 5865 19383 5899
rect 21005 5865 21039 5899
rect 21833 5865 21867 5899
rect 22017 5865 22051 5899
rect 2605 5797 2639 5831
rect 8769 5797 8803 5831
rect 10701 5797 10735 5831
rect 12173 5797 12207 5831
rect 14105 5797 14139 5831
rect 14289 5797 14323 5831
rect 18153 5797 18187 5831
rect 19533 5797 19567 5831
rect 18705 5729 18739 5763
rect 20269 5729 20303 5763
rect 20913 5729 20947 5763
rect 21557 5729 21591 5763
rect 1593 5661 1627 5695
rect 1869 5661 1903 5695
rect 2145 5661 2179 5695
rect 2513 5661 2547 5695
rect 2789 5661 2823 5695
rect 3249 5661 3283 5695
rect 3433 5661 3467 5695
rect 3985 5661 4019 5695
rect 4101 5663 4135 5697
rect 4353 5661 4387 5695
rect 6949 5661 6983 5695
rect 7205 5661 7239 5695
rect 7389 5661 7423 5695
rect 9229 5661 9263 5695
rect 9321 5661 9355 5695
rect 10793 5661 10827 5695
rect 11060 5661 11094 5695
rect 13737 5661 13771 5695
rect 14841 5661 14875 5695
rect 15025 5661 15059 5695
rect 16681 5661 16715 5695
rect 19073 5661 19107 5695
rect 19257 5661 19291 5695
rect 20177 5661 20211 5695
rect 21925 5661 21959 5695
rect 22569 5661 22603 5695
rect 22845 5661 22879 5695
rect 23305 5661 23339 5695
rect 1961 5593 1995 5627
rect 3525 5593 3559 5627
rect 4598 5593 4632 5627
rect 7634 5593 7668 5627
rect 9588 5593 9622 5627
rect 13470 5593 13504 5627
rect 14565 5593 14599 5627
rect 15292 5593 15326 5627
rect 16948 5593 16982 5627
rect 1777 5525 1811 5559
rect 3065 5525 3099 5559
rect 5733 5525 5767 5559
rect 5825 5525 5859 5559
rect 12357 5525 12391 5559
rect 16405 5525 16439 5559
rect 18061 5525 18095 5559
rect 2053 5321 2087 5355
rect 3157 5321 3191 5355
rect 5733 5321 5767 5355
rect 6101 5321 6135 5355
rect 14657 5321 14691 5355
rect 15117 5321 15151 5355
rect 15669 5321 15703 5355
rect 16313 5321 16347 5355
rect 17417 5321 17451 5355
rect 18797 5321 18831 5355
rect 21373 5321 21407 5355
rect 22201 5321 22235 5355
rect 23397 5321 23431 5355
rect 4169 5253 4203 5287
rect 6622 5253 6656 5287
rect 8576 5253 8610 5287
rect 11078 5253 11112 5287
rect 14933 5253 14967 5287
rect 1961 5185 1995 5219
rect 3341 5185 3375 5219
rect 4077 5185 4111 5219
rect 4609 5185 4643 5219
rect 6009 5185 6043 5219
rect 6377 5185 6411 5219
rect 13470 5185 13504 5219
rect 14381 5185 14415 5219
rect 14749 5185 14783 5219
rect 14841 5185 14875 5219
rect 15301 5185 15335 5219
rect 15761 5185 15795 5219
rect 16405 5185 16439 5219
rect 17233 5185 17267 5219
rect 18153 5185 18187 5219
rect 18889 5185 18923 5219
rect 21465 5185 21499 5219
rect 22753 5185 22787 5219
rect 23305 5185 23339 5219
rect 4353 5117 4387 5151
rect 8309 5117 8343 5151
rect 11345 5117 11379 5151
rect 13737 5117 13771 5151
rect 16681 5117 16715 5151
rect 18061 5117 18095 5151
rect 12357 5049 12391 5083
rect 18337 5049 18371 5083
rect 7757 4981 7791 5015
rect 9689 4981 9723 5015
rect 9965 4981 9999 5015
rect 13829 4981 13863 5015
rect 5825 4777 5859 4811
rect 6101 4777 6135 4811
rect 11253 4777 11287 4811
rect 13093 4777 13127 4811
rect 14289 4777 14323 4811
rect 16865 4777 16899 4811
rect 21741 4777 21775 4811
rect 22845 4777 22879 4811
rect 6469 4709 6503 4743
rect 9413 4709 9447 4743
rect 9505 4641 9539 4675
rect 12909 4641 12943 4675
rect 13369 4641 13403 4675
rect 22293 4641 22327 4675
rect 23489 4641 23523 4675
rect 5917 4573 5951 4607
rect 6009 4573 6043 4607
rect 6377 4573 6411 4607
rect 6653 4573 6687 4607
rect 7297 4573 7331 4607
rect 7389 4573 7423 4607
rect 7941 4573 7975 4607
rect 8677 4573 8711 4607
rect 9045 4573 9079 4607
rect 10977 4573 11011 4607
rect 11437 4573 11471 4607
rect 12653 4573 12687 4607
rect 13185 4573 13219 4607
rect 13461 4573 13495 4607
rect 14473 4573 14507 4607
rect 16957 4573 16991 4607
rect 10710 4505 10744 4539
rect 8125 4437 8159 4471
rect 9597 4437 9631 4471
rect 11529 4437 11563 4471
rect 9597 4233 9631 4267
rect 13093 4233 13127 4267
rect 12642 4165 12676 4199
rect 6469 4097 6503 4131
rect 6561 4097 6595 4131
rect 7113 4097 7147 4131
rect 8401 4097 8435 4131
rect 8861 4097 8895 4131
rect 9689 4097 9723 4131
rect 10241 4097 10275 4131
rect 10425 4097 10459 4131
rect 10517 4097 10551 4131
rect 11345 4097 11379 4131
rect 13185 4087 13219 4121
rect 22569 4097 22603 4131
rect 23213 4097 23247 4131
rect 7389 4029 7423 4063
rect 9045 4029 9079 4063
rect 10701 4029 10735 4063
rect 12909 4029 12943 4063
rect 8309 3961 8343 3995
rect 7297 3893 7331 3927
rect 8033 3893 8067 3927
rect 8677 3893 8711 3927
rect 11529 3893 11563 3927
rect 7573 3689 7607 3723
rect 8677 3689 8711 3723
rect 9045 3689 9079 3723
rect 10425 3689 10459 3723
rect 11897 3689 11931 3723
rect 12449 3689 12483 3723
rect 9137 3621 9171 3655
rect 9597 3621 9631 3655
rect 11529 3621 11563 3655
rect 12173 3553 12207 3587
rect 7665 3485 7699 3519
rect 8769 3485 8803 3519
rect 9505 3485 9539 3519
rect 10149 3485 10183 3519
rect 10517 3485 10551 3519
rect 11713 3485 11747 3519
rect 11989 3485 12023 3519
rect 12081 3485 12115 3519
rect 12541 3485 12575 3519
rect 11621 3009 11655 3043
rect 11897 2941 11931 2975
rect 7389 2465 7423 2499
rect 10701 2465 10735 2499
rect 7113 2397 7147 2431
rect 7941 2397 7975 2431
rect 10425 2397 10459 2431
rect 12541 2397 12575 2431
rect 13001 2397 13035 2431
rect 14197 2397 14231 2431
rect 17693 2397 17727 2431
rect 18245 2397 18279 2431
rect 8309 2329 8343 2363
rect 12173 2329 12207 2363
rect 13277 2329 13311 2363
rect 14565 2329 14599 2363
rect 17325 2329 17359 2363
rect 18613 2329 18647 2363
<< metal1 >>
rect 1104 24506 23828 24528
rect 1104 24454 1918 24506
rect 1970 24454 1982 24506
rect 2034 24454 2046 24506
rect 2098 24454 2110 24506
rect 2162 24454 2174 24506
rect 2226 24454 2238 24506
rect 2290 24454 7918 24506
rect 7970 24454 7982 24506
rect 8034 24454 8046 24506
rect 8098 24454 8110 24506
rect 8162 24454 8174 24506
rect 8226 24454 8238 24506
rect 8290 24454 13918 24506
rect 13970 24454 13982 24506
rect 14034 24454 14046 24506
rect 14098 24454 14110 24506
rect 14162 24454 14174 24506
rect 14226 24454 14238 24506
rect 14290 24454 19918 24506
rect 19970 24454 19982 24506
rect 20034 24454 20046 24506
rect 20098 24454 20110 24506
rect 20162 24454 20174 24506
rect 20226 24454 20238 24506
rect 20290 24454 23828 24506
rect 1104 24432 23828 24454
rect 7742 24216 7748 24268
rect 7800 24256 7806 24268
rect 8021 24259 8079 24265
rect 8021 24256 8033 24259
rect 7800 24228 8033 24256
rect 7800 24216 7806 24228
rect 8021 24225 8033 24228
rect 8067 24225 8079 24259
rect 8021 24219 8079 24225
rect 8386 24216 8392 24268
rect 8444 24256 8450 24268
rect 9309 24259 9367 24265
rect 9309 24256 9321 24259
rect 8444 24228 9321 24256
rect 8444 24216 8450 24228
rect 9309 24225 9321 24228
rect 9355 24225 9367 24259
rect 9309 24219 9367 24225
rect 10962 24216 10968 24268
rect 11020 24256 11026 24268
rect 11885 24259 11943 24265
rect 11885 24256 11897 24259
rect 11020 24228 11897 24256
rect 11020 24216 11026 24228
rect 11885 24225 11897 24228
rect 11931 24225 11943 24259
rect 11885 24219 11943 24225
rect 13538 24216 13544 24268
rect 13596 24256 13602 24268
rect 14277 24259 14335 24265
rect 14277 24256 14289 24259
rect 13596 24228 14289 24256
rect 13596 24216 13602 24228
rect 14277 24225 14289 24228
rect 14323 24225 14335 24259
rect 14277 24219 14335 24225
rect 14458 24216 14464 24268
rect 14516 24256 14522 24268
rect 14516 24228 14780 24256
rect 14516 24216 14522 24228
rect 7558 24148 7564 24200
rect 7616 24188 7622 24200
rect 7837 24191 7895 24197
rect 7837 24188 7849 24191
rect 7616 24160 7849 24188
rect 7616 24148 7622 24160
rect 7837 24157 7849 24160
rect 7883 24157 7895 24191
rect 7837 24151 7895 24157
rect 9033 24191 9091 24197
rect 9033 24157 9045 24191
rect 9079 24188 9091 24191
rect 9582 24188 9588 24200
rect 9079 24160 9588 24188
rect 9079 24157 9091 24160
rect 9033 24151 9091 24157
rect 9582 24148 9588 24160
rect 9640 24148 9646 24200
rect 10778 24148 10784 24200
rect 10836 24188 10842 24200
rect 11609 24191 11667 24197
rect 11609 24188 11621 24191
rect 10836 24160 11621 24188
rect 10836 24148 10842 24160
rect 11609 24157 11621 24160
rect 11655 24157 11667 24191
rect 11609 24151 11667 24157
rect 12986 24148 12992 24200
rect 13044 24188 13050 24200
rect 14093 24191 14151 24197
rect 14093 24188 14105 24191
rect 13044 24160 14105 24188
rect 13044 24148 13050 24160
rect 14093 24157 14105 24160
rect 14139 24157 14151 24191
rect 14093 24151 14151 24157
rect 14550 24148 14556 24200
rect 14608 24188 14614 24200
rect 14645 24191 14703 24197
rect 14645 24188 14657 24191
rect 14608 24160 14657 24188
rect 14608 24148 14614 24160
rect 14645 24157 14657 24160
rect 14691 24157 14703 24191
rect 14752 24188 14780 24228
rect 14826 24216 14832 24268
rect 14884 24256 14890 24268
rect 15565 24259 15623 24265
rect 15565 24256 15577 24259
rect 14884 24228 15577 24256
rect 14884 24216 14890 24228
rect 15565 24225 15577 24228
rect 15611 24225 15623 24259
rect 15565 24219 15623 24225
rect 14921 24191 14979 24197
rect 14921 24188 14933 24191
rect 14752 24160 14933 24188
rect 14645 24151 14703 24157
rect 14921 24157 14933 24160
rect 14967 24157 14979 24191
rect 14921 24151 14979 24157
rect 15289 24191 15347 24197
rect 15289 24157 15301 24191
rect 15335 24188 15347 24191
rect 15378 24188 15384 24200
rect 15335 24160 15384 24188
rect 15335 24157 15347 24160
rect 15289 24151 15347 24157
rect 15378 24148 15384 24160
rect 15436 24148 15442 24200
rect 1104 23962 23828 23984
rect 1104 23910 2658 23962
rect 2710 23910 2722 23962
rect 2774 23910 2786 23962
rect 2838 23910 2850 23962
rect 2902 23910 2914 23962
rect 2966 23910 2978 23962
rect 3030 23910 8658 23962
rect 8710 23910 8722 23962
rect 8774 23910 8786 23962
rect 8838 23910 8850 23962
rect 8902 23910 8914 23962
rect 8966 23910 8978 23962
rect 9030 23910 14658 23962
rect 14710 23910 14722 23962
rect 14774 23910 14786 23962
rect 14838 23910 14850 23962
rect 14902 23910 14914 23962
rect 14966 23910 14978 23962
rect 15030 23910 20658 23962
rect 20710 23910 20722 23962
rect 20774 23910 20786 23962
rect 20838 23910 20850 23962
rect 20902 23910 20914 23962
rect 20966 23910 20978 23962
rect 21030 23910 23828 23962
rect 1104 23888 23828 23910
rect 1104 23418 23828 23440
rect 1104 23366 1918 23418
rect 1970 23366 1982 23418
rect 2034 23366 2046 23418
rect 2098 23366 2110 23418
rect 2162 23366 2174 23418
rect 2226 23366 2238 23418
rect 2290 23366 7918 23418
rect 7970 23366 7982 23418
rect 8034 23366 8046 23418
rect 8098 23366 8110 23418
rect 8162 23366 8174 23418
rect 8226 23366 8238 23418
rect 8290 23366 13918 23418
rect 13970 23366 13982 23418
rect 14034 23366 14046 23418
rect 14098 23366 14110 23418
rect 14162 23366 14174 23418
rect 14226 23366 14238 23418
rect 14290 23366 19918 23418
rect 19970 23366 19982 23418
rect 20034 23366 20046 23418
rect 20098 23366 20110 23418
rect 20162 23366 20174 23418
rect 20226 23366 20238 23418
rect 20290 23366 23828 23418
rect 1104 23344 23828 23366
rect 1104 22874 23828 22896
rect 1104 22822 2658 22874
rect 2710 22822 2722 22874
rect 2774 22822 2786 22874
rect 2838 22822 2850 22874
rect 2902 22822 2914 22874
rect 2966 22822 2978 22874
rect 3030 22822 8658 22874
rect 8710 22822 8722 22874
rect 8774 22822 8786 22874
rect 8838 22822 8850 22874
rect 8902 22822 8914 22874
rect 8966 22822 8978 22874
rect 9030 22822 14658 22874
rect 14710 22822 14722 22874
rect 14774 22822 14786 22874
rect 14838 22822 14850 22874
rect 14902 22822 14914 22874
rect 14966 22822 14978 22874
rect 15030 22822 20658 22874
rect 20710 22822 20722 22874
rect 20774 22822 20786 22874
rect 20838 22822 20850 22874
rect 20902 22822 20914 22874
rect 20966 22822 20978 22874
rect 21030 22822 23828 22874
rect 1104 22800 23828 22822
rect 11241 22627 11299 22633
rect 11241 22593 11253 22627
rect 11287 22624 11299 22627
rect 16482 22624 16488 22636
rect 11287 22596 16488 22624
rect 11287 22593 11299 22596
rect 11241 22587 11299 22593
rect 16482 22584 16488 22596
rect 16540 22584 16546 22636
rect 10962 22380 10968 22432
rect 11020 22420 11026 22432
rect 11057 22423 11115 22429
rect 11057 22420 11069 22423
rect 11020 22392 11069 22420
rect 11020 22380 11026 22392
rect 11057 22389 11069 22392
rect 11103 22389 11115 22423
rect 11057 22383 11115 22389
rect 1104 22330 23828 22352
rect 1104 22278 1918 22330
rect 1970 22278 1982 22330
rect 2034 22278 2046 22330
rect 2098 22278 2110 22330
rect 2162 22278 2174 22330
rect 2226 22278 2238 22330
rect 2290 22278 7918 22330
rect 7970 22278 7982 22330
rect 8034 22278 8046 22330
rect 8098 22278 8110 22330
rect 8162 22278 8174 22330
rect 8226 22278 8238 22330
rect 8290 22278 13918 22330
rect 13970 22278 13982 22330
rect 14034 22278 14046 22330
rect 14098 22278 14110 22330
rect 14162 22278 14174 22330
rect 14226 22278 14238 22330
rect 14290 22278 19918 22330
rect 19970 22278 19982 22330
rect 20034 22278 20046 22330
rect 20098 22278 20110 22330
rect 20162 22278 20174 22330
rect 20226 22278 20238 22330
rect 20290 22278 23828 22330
rect 1104 22256 23828 22278
rect 9861 22151 9919 22157
rect 9861 22117 9873 22151
rect 9907 22148 9919 22151
rect 10318 22148 10324 22160
rect 9907 22120 10324 22148
rect 9907 22117 9919 22120
rect 9861 22111 9919 22117
rect 10318 22108 10324 22120
rect 10376 22108 10382 22160
rect 9677 22083 9735 22089
rect 9677 22049 9689 22083
rect 9723 22080 9735 22083
rect 10042 22080 10048 22092
rect 9723 22052 10048 22080
rect 9723 22049 9735 22052
rect 9677 22043 9735 22049
rect 10042 22040 10048 22052
rect 10100 22040 10106 22092
rect 8481 22015 8539 22021
rect 8481 22012 8493 22015
rect 7852 21984 8493 22012
rect 7852 21956 7880 21984
rect 8481 21981 8493 21984
rect 8527 21981 8539 22015
rect 8481 21975 8539 21981
rect 8757 22015 8815 22021
rect 8757 21981 8769 22015
rect 8803 22012 8815 22015
rect 8803 21984 9904 22012
rect 8803 21981 8815 21984
rect 8757 21975 8815 21981
rect 7834 21904 7840 21956
rect 7892 21904 7898 21956
rect 6822 21836 6828 21888
rect 6880 21876 6886 21888
rect 8389 21879 8447 21885
rect 8389 21876 8401 21879
rect 6880 21848 8401 21876
rect 6880 21836 6886 21848
rect 8389 21845 8401 21848
rect 8435 21845 8447 21879
rect 8389 21839 8447 21845
rect 8570 21836 8576 21888
rect 8628 21876 8634 21888
rect 8665 21879 8723 21885
rect 8665 21876 8677 21879
rect 8628 21848 8677 21876
rect 8628 21836 8634 21848
rect 8665 21845 8677 21848
rect 8711 21845 8723 21879
rect 9876 21876 9904 21984
rect 9950 21972 9956 22024
rect 10008 22012 10014 22024
rect 10689 22015 10747 22021
rect 10689 22012 10701 22015
rect 10008 21984 10701 22012
rect 10008 21972 10014 21984
rect 10689 21981 10701 21984
rect 10735 21981 10747 22015
rect 12345 22015 12403 22021
rect 10689 21975 10747 21981
rect 10888 21984 12112 22012
rect 10137 21947 10195 21953
rect 10137 21913 10149 21947
rect 10183 21944 10195 21947
rect 10502 21944 10508 21956
rect 10183 21916 10508 21944
rect 10183 21913 10195 21916
rect 10137 21907 10195 21913
rect 10502 21904 10508 21916
rect 10560 21904 10566 21956
rect 10594 21904 10600 21956
rect 10652 21944 10658 21956
rect 10888 21944 10916 21984
rect 10962 21953 10968 21956
rect 10652 21916 10916 21944
rect 10652 21904 10658 21916
rect 10956 21907 10968 21953
rect 10962 21904 10968 21907
rect 11020 21904 11026 21956
rect 12084 21944 12112 21984
rect 12345 21981 12357 22015
rect 12391 21981 12403 22015
rect 12345 21975 12403 21981
rect 12360 21944 12388 21975
rect 12618 21972 12624 22024
rect 12676 21972 12682 22024
rect 14274 21972 14280 22024
rect 14332 21972 14338 22024
rect 14369 22015 14427 22021
rect 14369 21981 14381 22015
rect 14415 21981 14427 22015
rect 14369 21975 14427 21981
rect 15197 22015 15255 22021
rect 15197 21981 15209 22015
rect 15243 22012 15255 22015
rect 15243 21984 15516 22012
rect 15243 21981 15255 21984
rect 15197 21975 15255 21981
rect 13170 21944 13176 21956
rect 12084 21916 12204 21944
rect 12360 21916 13176 21944
rect 11054 21876 11060 21888
rect 9876 21848 11060 21876
rect 8665 21839 8723 21845
rect 11054 21836 11060 21848
rect 11112 21836 11118 21888
rect 12066 21836 12072 21888
rect 12124 21836 12130 21888
rect 12176 21885 12204 21916
rect 13170 21904 13176 21916
rect 13228 21904 13234 21956
rect 14384 21944 14412 21975
rect 13740 21916 14412 21944
rect 13740 21888 13768 21916
rect 15488 21888 15516 21984
rect 12161 21879 12219 21885
rect 12161 21845 12173 21879
rect 12207 21845 12219 21879
rect 12161 21839 12219 21845
rect 13262 21836 13268 21888
rect 13320 21836 13326 21888
rect 13722 21836 13728 21888
rect 13780 21836 13786 21888
rect 13814 21836 13820 21888
rect 13872 21876 13878 21888
rect 14185 21879 14243 21885
rect 14185 21876 14197 21879
rect 13872 21848 14197 21876
rect 13872 21836 13878 21848
rect 14185 21845 14197 21848
rect 14231 21845 14243 21879
rect 14185 21839 14243 21845
rect 14458 21836 14464 21888
rect 14516 21836 14522 21888
rect 15286 21836 15292 21888
rect 15344 21836 15350 21888
rect 15470 21836 15476 21888
rect 15528 21836 15534 21888
rect 1104 21786 23828 21808
rect 1104 21734 2658 21786
rect 2710 21734 2722 21786
rect 2774 21734 2786 21786
rect 2838 21734 2850 21786
rect 2902 21734 2914 21786
rect 2966 21734 2978 21786
rect 3030 21734 8658 21786
rect 8710 21734 8722 21786
rect 8774 21734 8786 21786
rect 8838 21734 8850 21786
rect 8902 21734 8914 21786
rect 8966 21734 8978 21786
rect 9030 21734 14658 21786
rect 14710 21734 14722 21786
rect 14774 21734 14786 21786
rect 14838 21734 14850 21786
rect 14902 21734 14914 21786
rect 14966 21734 14978 21786
rect 15030 21734 20658 21786
rect 20710 21734 20722 21786
rect 20774 21734 20786 21786
rect 20838 21734 20850 21786
rect 20902 21734 20914 21786
rect 20966 21734 20978 21786
rect 21030 21734 23828 21786
rect 1104 21712 23828 21734
rect 10318 21632 10324 21684
rect 10376 21632 10382 21684
rect 10502 21632 10508 21684
rect 10560 21672 10566 21684
rect 11882 21672 11888 21684
rect 10560 21644 11888 21672
rect 10560 21632 10566 21644
rect 11882 21632 11888 21644
rect 11940 21632 11946 21684
rect 11054 21564 11060 21616
rect 11112 21604 11118 21616
rect 13722 21604 13728 21616
rect 11112 21576 13728 21604
rect 11112 21564 11118 21576
rect 13722 21564 13728 21576
rect 13780 21604 13786 21616
rect 13780 21576 14412 21604
rect 13780 21564 13786 21576
rect 5626 21496 5632 21548
rect 5684 21536 5690 21548
rect 6805 21539 6863 21545
rect 6805 21536 6817 21539
rect 5684 21508 6817 21536
rect 5684 21496 5690 21508
rect 6805 21505 6817 21508
rect 6851 21505 6863 21539
rect 6805 21499 6863 21505
rect 10502 21496 10508 21548
rect 10560 21536 10566 21548
rect 11149 21539 11207 21545
rect 11149 21536 11161 21539
rect 10560 21508 11161 21536
rect 10560 21496 10566 21508
rect 11149 21505 11161 21508
rect 11195 21505 11207 21539
rect 11149 21499 11207 21505
rect 11517 21539 11575 21545
rect 11517 21505 11529 21539
rect 11563 21505 11575 21539
rect 11517 21499 11575 21505
rect 6546 21428 6552 21480
rect 6604 21428 6610 21480
rect 7650 21428 7656 21480
rect 7708 21468 7714 21480
rect 8021 21471 8079 21477
rect 8021 21468 8033 21471
rect 7708 21440 8033 21468
rect 7708 21428 7714 21440
rect 8021 21437 8033 21440
rect 8067 21437 8079 21471
rect 8021 21431 8079 21437
rect 9401 21471 9459 21477
rect 9401 21437 9413 21471
rect 9447 21468 9459 21471
rect 9490 21468 9496 21480
rect 9447 21440 9496 21468
rect 9447 21437 9459 21440
rect 9401 21431 9459 21437
rect 9490 21428 9496 21440
rect 9548 21428 9554 21480
rect 9766 21428 9772 21480
rect 9824 21428 9830 21480
rect 10410 21428 10416 21480
rect 10468 21428 10474 21480
rect 11532 21400 11560 21499
rect 11606 21496 11612 21548
rect 11664 21536 11670 21548
rect 12529 21539 12587 21545
rect 12529 21536 12541 21539
rect 11664 21508 12541 21536
rect 11664 21496 11670 21508
rect 12529 21505 12541 21508
rect 12575 21505 12587 21539
rect 12529 21499 12587 21505
rect 12618 21496 12624 21548
rect 12676 21536 12682 21548
rect 14384 21545 14412 21576
rect 12785 21539 12843 21545
rect 12785 21536 12797 21539
rect 12676 21508 12797 21536
rect 12676 21496 12682 21508
rect 12785 21505 12797 21508
rect 12831 21505 12843 21539
rect 12785 21499 12843 21505
rect 14369 21539 14427 21545
rect 14369 21505 14381 21539
rect 14415 21505 14427 21539
rect 14369 21499 14427 21505
rect 15470 21496 15476 21548
rect 15528 21496 15534 21548
rect 11790 21428 11796 21480
rect 11848 21428 11854 21480
rect 14550 21428 14556 21480
rect 14608 21428 14614 21480
rect 15562 21428 15568 21480
rect 15620 21468 15626 21480
rect 15657 21471 15715 21477
rect 15657 21468 15669 21471
rect 15620 21440 15669 21468
rect 15620 21428 15626 21440
rect 15657 21437 15669 21440
rect 15703 21437 15715 21471
rect 15657 21431 15715 21437
rect 17218 21428 17224 21480
rect 17276 21428 17282 21480
rect 18138 21428 18144 21480
rect 18196 21428 18202 21480
rect 9416 21372 11560 21400
rect 9416 21344 9444 21372
rect 7742 21292 7748 21344
rect 7800 21332 7806 21344
rect 7929 21335 7987 21341
rect 7929 21332 7941 21335
rect 7800 21304 7941 21332
rect 7800 21292 7806 21304
rect 7929 21301 7941 21304
rect 7975 21301 7987 21335
rect 7929 21295 7987 21301
rect 8478 21292 8484 21344
rect 8536 21332 8542 21344
rect 8665 21335 8723 21341
rect 8665 21332 8677 21335
rect 8536 21304 8677 21332
rect 8536 21292 8542 21304
rect 8665 21301 8677 21304
rect 8711 21301 8723 21335
rect 8665 21295 8723 21301
rect 8757 21335 8815 21341
rect 8757 21301 8769 21335
rect 8803 21332 8815 21335
rect 9306 21332 9312 21344
rect 8803 21304 9312 21332
rect 8803 21301 8815 21304
rect 8757 21295 8815 21301
rect 9306 21292 9312 21304
rect 9364 21292 9370 21344
rect 9398 21292 9404 21344
rect 9456 21292 9462 21344
rect 11057 21335 11115 21341
rect 11057 21301 11069 21335
rect 11103 21332 11115 21335
rect 11146 21332 11152 21344
rect 11103 21304 11152 21332
rect 11103 21301 11115 21304
rect 11057 21295 11115 21301
rect 11146 21292 11152 21304
rect 11204 21292 11210 21344
rect 11238 21292 11244 21344
rect 11296 21292 11302 21344
rect 11606 21292 11612 21344
rect 11664 21292 11670 21344
rect 12434 21292 12440 21344
rect 12492 21292 12498 21344
rect 13722 21292 13728 21344
rect 13780 21332 13786 21344
rect 13909 21335 13967 21341
rect 13909 21332 13921 21335
rect 13780 21304 13921 21332
rect 13780 21292 13786 21304
rect 13909 21301 13921 21304
rect 13955 21301 13967 21335
rect 13909 21295 13967 21301
rect 14277 21335 14335 21341
rect 14277 21301 14289 21335
rect 14323 21332 14335 21335
rect 14734 21332 14740 21344
rect 14323 21304 14740 21332
rect 14323 21301 14335 21304
rect 14277 21295 14335 21301
rect 14734 21292 14740 21304
rect 14792 21292 14798 21344
rect 15194 21292 15200 21344
rect 15252 21292 15258 21344
rect 15378 21292 15384 21344
rect 15436 21292 15442 21344
rect 16298 21292 16304 21344
rect 16356 21292 16362 21344
rect 16666 21292 16672 21344
rect 16724 21292 16730 21344
rect 18782 21292 18788 21344
rect 18840 21292 18846 21344
rect 1104 21242 23828 21264
rect 1104 21190 1918 21242
rect 1970 21190 1982 21242
rect 2034 21190 2046 21242
rect 2098 21190 2110 21242
rect 2162 21190 2174 21242
rect 2226 21190 2238 21242
rect 2290 21190 7918 21242
rect 7970 21190 7982 21242
rect 8034 21190 8046 21242
rect 8098 21190 8110 21242
rect 8162 21190 8174 21242
rect 8226 21190 8238 21242
rect 8290 21190 13918 21242
rect 13970 21190 13982 21242
rect 14034 21190 14046 21242
rect 14098 21190 14110 21242
rect 14162 21190 14174 21242
rect 14226 21190 14238 21242
rect 14290 21190 19918 21242
rect 19970 21190 19982 21242
rect 20034 21190 20046 21242
rect 20098 21190 20110 21242
rect 20162 21190 20174 21242
rect 20226 21190 20238 21242
rect 20290 21190 23828 21242
rect 1104 21168 23828 21190
rect 10962 21088 10968 21140
rect 11020 21088 11026 21140
rect 11238 21128 11244 21140
rect 11072 21100 11244 21128
rect 5534 20952 5540 21004
rect 5592 20992 5598 21004
rect 6178 20992 6184 21004
rect 5592 20964 6184 20992
rect 5592 20952 5598 20964
rect 6178 20952 6184 20964
rect 6236 20992 6242 21004
rect 6546 20992 6552 21004
rect 6236 20964 6552 20992
rect 6236 20952 6242 20964
rect 6546 20952 6552 20964
rect 6604 20992 6610 21004
rect 11072 21001 11100 21100
rect 11238 21088 11244 21100
rect 11296 21088 11302 21140
rect 12434 21088 12440 21140
rect 12492 21088 12498 21140
rect 14734 21128 14740 21140
rect 14108 21100 14740 21128
rect 6825 20995 6883 21001
rect 6825 20992 6837 20995
rect 6604 20964 6837 20992
rect 6604 20952 6610 20964
rect 6825 20961 6837 20964
rect 6871 20961 6883 20995
rect 11057 20995 11115 21001
rect 6825 20955 6883 20961
rect 8220 20964 8616 20992
rect 4249 20927 4307 20933
rect 4249 20893 4261 20927
rect 4295 20893 4307 20927
rect 4249 20887 4307 20893
rect 4341 20927 4399 20933
rect 4341 20893 4353 20927
rect 4387 20924 4399 20927
rect 4525 20927 4583 20933
rect 4525 20924 4537 20927
rect 4387 20896 4537 20924
rect 4387 20893 4399 20896
rect 4341 20887 4399 20893
rect 4525 20893 4537 20896
rect 4571 20893 4583 20927
rect 4525 20887 4583 20893
rect 6089 20927 6147 20933
rect 6089 20893 6101 20927
rect 6135 20924 6147 20927
rect 6730 20924 6736 20936
rect 6135 20896 6736 20924
rect 6135 20893 6147 20896
rect 6089 20887 6147 20893
rect 4264 20856 4292 20887
rect 6730 20884 6736 20896
rect 6788 20924 6794 20936
rect 7081 20927 7139 20933
rect 7081 20924 7093 20927
rect 6788 20896 7093 20924
rect 6788 20884 6794 20896
rect 7081 20893 7093 20896
rect 7127 20893 7139 20927
rect 7834 20924 7840 20936
rect 7081 20887 7139 20893
rect 7208 20896 7840 20924
rect 4792 20859 4850 20865
rect 4264 20828 4384 20856
rect 4356 20800 4384 20828
rect 4792 20825 4804 20859
rect 4838 20856 4850 20859
rect 4890 20856 4896 20868
rect 4838 20828 4896 20856
rect 4838 20825 4850 20828
rect 4792 20819 4850 20825
rect 4890 20816 4896 20828
rect 4948 20816 4954 20868
rect 7208 20856 7236 20896
rect 7834 20884 7840 20896
rect 7892 20924 7898 20936
rect 8220 20924 8248 20964
rect 8588 20933 8616 20964
rect 9140 20964 9720 20992
rect 9140 20933 9168 20964
rect 8481 20927 8539 20933
rect 8481 20924 8493 20927
rect 7892 20896 8248 20924
rect 8312 20896 8493 20924
rect 7892 20884 7898 20896
rect 7024 20828 7236 20856
rect 7024 20800 7052 20828
rect 8312 20800 8340 20896
rect 8481 20893 8493 20896
rect 8527 20893 8539 20927
rect 8481 20887 8539 20893
rect 8573 20927 8631 20933
rect 8573 20893 8585 20927
rect 8619 20893 8631 20927
rect 8573 20887 8631 20893
rect 9125 20927 9183 20933
rect 9125 20893 9137 20927
rect 9171 20893 9183 20927
rect 9125 20887 9183 20893
rect 9309 20927 9367 20933
rect 9309 20893 9321 20927
rect 9355 20893 9367 20927
rect 9309 20887 9367 20893
rect 9401 20927 9459 20933
rect 9401 20893 9413 20927
rect 9447 20924 9459 20927
rect 9585 20927 9643 20933
rect 9585 20924 9597 20927
rect 9447 20896 9597 20924
rect 9447 20893 9459 20896
rect 9401 20887 9459 20893
rect 9585 20893 9597 20896
rect 9631 20893 9643 20927
rect 9692 20924 9720 20964
rect 11057 20961 11069 20995
rect 11103 20961 11115 20995
rect 12452 20992 12480 21088
rect 14108 21001 14136 21100
rect 14734 21088 14740 21100
rect 14792 21088 14798 21140
rect 15286 21088 15292 21140
rect 15344 21088 15350 21140
rect 15473 21131 15531 21137
rect 15473 21097 15485 21131
rect 15519 21128 15531 21131
rect 15562 21128 15568 21140
rect 15519 21100 15568 21128
rect 15519 21097 15531 21100
rect 15473 21091 15531 21097
rect 15562 21088 15568 21100
rect 15620 21088 15626 21140
rect 14093 20995 14151 21001
rect 12452 20964 12664 20992
rect 11057 20955 11115 20961
rect 9692 20896 11100 20924
rect 9585 20887 9643 20893
rect 8665 20859 8723 20865
rect 8665 20825 8677 20859
rect 8711 20856 8723 20859
rect 9214 20856 9220 20868
rect 8711 20828 9220 20856
rect 8711 20825 8723 20828
rect 8665 20819 8723 20825
rect 9214 20816 9220 20828
rect 9272 20816 9278 20868
rect 9324 20856 9352 20887
rect 9852 20859 9910 20865
rect 9324 20828 9444 20856
rect 9416 20800 9444 20828
rect 9852 20825 9864 20859
rect 9898 20856 9910 20859
rect 10594 20856 10600 20868
rect 9898 20828 10600 20856
rect 9898 20825 9910 20828
rect 9852 20819 9910 20825
rect 10594 20816 10600 20828
rect 10652 20816 10658 20868
rect 11072 20800 11100 20896
rect 12526 20884 12532 20936
rect 12584 20884 12590 20936
rect 12636 20924 12664 20964
rect 14093 20961 14105 20995
rect 14139 20961 14151 20995
rect 15304 20992 15332 21088
rect 16945 21063 17003 21069
rect 16945 21029 16957 21063
rect 16991 21029 17003 21063
rect 16945 21023 17003 21029
rect 15565 20995 15623 21001
rect 15565 20992 15577 20995
rect 15304 20964 15577 20992
rect 14093 20955 14151 20961
rect 15565 20961 15577 20964
rect 15611 20961 15623 20995
rect 16960 20992 16988 21023
rect 17589 20995 17647 21001
rect 17589 20992 17601 20995
rect 16960 20964 17601 20992
rect 15565 20955 15623 20961
rect 17589 20961 17601 20964
rect 17635 20961 17647 20995
rect 17589 20955 17647 20961
rect 17972 20964 19288 20992
rect 12785 20927 12843 20933
rect 12785 20924 12797 20927
rect 12636 20896 12797 20924
rect 12785 20893 12797 20896
rect 12831 20893 12843 20927
rect 12785 20887 12843 20893
rect 13722 20884 13728 20936
rect 13780 20924 13786 20936
rect 14349 20927 14407 20933
rect 14349 20924 14361 20927
rect 13780 20896 14361 20924
rect 13780 20884 13786 20896
rect 14349 20893 14361 20896
rect 14395 20893 14407 20927
rect 14349 20887 14407 20893
rect 14642 20884 14648 20936
rect 14700 20884 14706 20936
rect 15832 20927 15890 20933
rect 15832 20893 15844 20927
rect 15878 20924 15890 20927
rect 16298 20924 16304 20936
rect 15878 20896 16304 20924
rect 15878 20893 15890 20896
rect 15832 20887 15890 20893
rect 16298 20884 16304 20896
rect 16356 20884 16362 20936
rect 17770 20884 17776 20936
rect 17828 20924 17834 20936
rect 17972 20933 18000 20964
rect 17957 20927 18015 20933
rect 17957 20924 17969 20927
rect 17828 20896 17969 20924
rect 17828 20884 17834 20896
rect 17957 20893 17969 20896
rect 18003 20893 18015 20927
rect 17957 20887 18015 20893
rect 18325 20927 18383 20933
rect 18325 20893 18337 20927
rect 18371 20924 18383 20927
rect 18414 20924 18420 20936
rect 18371 20896 18420 20924
rect 18371 20893 18383 20896
rect 18325 20887 18383 20893
rect 18414 20884 18420 20896
rect 18472 20884 18478 20936
rect 19260 20933 19288 20964
rect 19245 20927 19303 20933
rect 19245 20893 19257 20927
rect 19291 20893 19303 20927
rect 19245 20887 19303 20893
rect 11330 20865 11336 20868
rect 11324 20819 11336 20865
rect 11330 20816 11336 20819
rect 11388 20816 11394 20868
rect 4338 20748 4344 20800
rect 4396 20748 4402 20800
rect 5350 20748 5356 20800
rect 5408 20788 5414 20800
rect 5905 20791 5963 20797
rect 5905 20788 5917 20791
rect 5408 20760 5917 20788
rect 5408 20748 5414 20760
rect 5905 20757 5917 20760
rect 5951 20757 5963 20791
rect 5905 20751 5963 20757
rect 6733 20791 6791 20797
rect 6733 20757 6745 20791
rect 6779 20788 6791 20791
rect 6914 20788 6920 20800
rect 6779 20760 6920 20788
rect 6779 20757 6791 20760
rect 6733 20751 6791 20757
rect 6914 20748 6920 20760
rect 6972 20748 6978 20800
rect 7006 20748 7012 20800
rect 7064 20748 7070 20800
rect 7834 20748 7840 20800
rect 7892 20788 7898 20800
rect 8205 20791 8263 20797
rect 8205 20788 8217 20791
rect 7892 20760 8217 20788
rect 7892 20748 7898 20760
rect 8205 20757 8217 20760
rect 8251 20757 8263 20791
rect 8205 20751 8263 20757
rect 8294 20748 8300 20800
rect 8352 20748 8358 20800
rect 8386 20748 8392 20800
rect 8444 20748 8450 20800
rect 9033 20791 9091 20797
rect 9033 20757 9045 20791
rect 9079 20788 9091 20791
rect 9122 20788 9128 20800
rect 9079 20760 9128 20788
rect 9079 20757 9091 20760
rect 9033 20751 9091 20757
rect 9122 20748 9128 20760
rect 9180 20748 9186 20800
rect 9398 20748 9404 20800
rect 9456 20748 9462 20800
rect 11054 20748 11060 20800
rect 11112 20748 11118 20800
rect 11790 20748 11796 20800
rect 11848 20788 11854 20800
rect 12437 20791 12495 20797
rect 12437 20788 12449 20791
rect 11848 20760 12449 20788
rect 11848 20748 11854 20760
rect 12437 20757 12449 20760
rect 12483 20757 12495 20791
rect 12437 20751 12495 20757
rect 13909 20791 13967 20797
rect 13909 20757 13921 20791
rect 13955 20788 13967 20791
rect 14660 20788 14688 20884
rect 18877 20859 18935 20865
rect 18877 20825 18889 20859
rect 18923 20856 18935 20859
rect 19518 20856 19524 20868
rect 18923 20828 19524 20856
rect 18923 20825 18935 20828
rect 18877 20819 18935 20825
rect 19518 20816 19524 20828
rect 19576 20816 19582 20868
rect 13955 20760 14688 20788
rect 13955 20757 13967 20760
rect 13909 20751 13967 20757
rect 15562 20748 15568 20800
rect 15620 20788 15626 20800
rect 17037 20791 17095 20797
rect 17037 20788 17049 20791
rect 15620 20760 17049 20788
rect 15620 20748 15626 20760
rect 17037 20757 17049 20760
rect 17083 20757 17095 20791
rect 17037 20751 17095 20757
rect 18046 20748 18052 20800
rect 18104 20748 18110 20800
rect 19334 20748 19340 20800
rect 19392 20748 19398 20800
rect 1104 20698 23828 20720
rect 1104 20646 2658 20698
rect 2710 20646 2722 20698
rect 2774 20646 2786 20698
rect 2838 20646 2850 20698
rect 2902 20646 2914 20698
rect 2966 20646 2978 20698
rect 3030 20646 8658 20698
rect 8710 20646 8722 20698
rect 8774 20646 8786 20698
rect 8838 20646 8850 20698
rect 8902 20646 8914 20698
rect 8966 20646 8978 20698
rect 9030 20646 14658 20698
rect 14710 20646 14722 20698
rect 14774 20646 14786 20698
rect 14838 20646 14850 20698
rect 14902 20646 14914 20698
rect 14966 20646 14978 20698
rect 15030 20646 20658 20698
rect 20710 20646 20722 20698
rect 20774 20646 20786 20698
rect 20838 20646 20850 20698
rect 20902 20646 20914 20698
rect 20966 20646 20978 20698
rect 21030 20646 23828 20698
rect 1104 20624 23828 20646
rect 8294 20584 8300 20596
rect 6748 20556 8300 20584
rect 4816 20488 5488 20516
rect 4816 20460 4844 20488
rect 5460 20460 5488 20488
rect 4798 20408 4804 20460
rect 4856 20408 4862 20460
rect 5068 20451 5126 20457
rect 5068 20417 5080 20451
rect 5114 20448 5126 20451
rect 5350 20448 5356 20460
rect 5114 20420 5356 20448
rect 5114 20417 5126 20420
rect 5068 20411 5126 20417
rect 5350 20408 5356 20420
rect 5408 20408 5414 20460
rect 5442 20408 5448 20460
rect 5500 20408 5506 20460
rect 6457 20451 6515 20457
rect 6457 20448 6469 20451
rect 6288 20420 6469 20448
rect 6288 20324 6316 20420
rect 6457 20417 6469 20420
rect 6503 20417 6515 20451
rect 6457 20411 6515 20417
rect 6638 20408 6644 20460
rect 6696 20448 6702 20460
rect 6748 20457 6776 20556
rect 8294 20544 8300 20556
rect 8352 20584 8358 20596
rect 8662 20584 8668 20596
rect 8352 20556 8668 20584
rect 8352 20544 8358 20556
rect 8662 20544 8668 20556
rect 8720 20544 8726 20596
rect 9861 20587 9919 20593
rect 9861 20553 9873 20587
rect 9907 20584 9919 20587
rect 10410 20584 10416 20596
rect 9907 20556 10416 20584
rect 9907 20553 9919 20556
rect 9861 20547 9919 20553
rect 10410 20544 10416 20556
rect 10468 20544 10474 20596
rect 11330 20544 11336 20596
rect 11388 20544 11394 20596
rect 14458 20584 14464 20596
rect 13004 20556 14464 20584
rect 6825 20519 6883 20525
rect 6825 20485 6837 20519
rect 6871 20516 6883 20519
rect 8748 20519 8806 20525
rect 6871 20488 8524 20516
rect 6871 20485 6883 20488
rect 6825 20479 6883 20485
rect 6733 20451 6791 20457
rect 6733 20448 6745 20451
rect 6696 20420 6745 20448
rect 6696 20408 6702 20420
rect 6733 20417 6745 20420
rect 6779 20417 6791 20451
rect 6733 20411 6791 20417
rect 7742 20408 7748 20460
rect 7800 20448 7806 20460
rect 8496 20457 8524 20488
rect 8748 20485 8760 20519
rect 8794 20516 8806 20519
rect 9306 20516 9312 20528
rect 8794 20488 9312 20516
rect 8794 20485 8806 20488
rect 8748 20479 8806 20485
rect 9306 20476 9312 20488
rect 9364 20476 9370 20528
rect 11790 20525 11796 20528
rect 11784 20516 11796 20525
rect 11751 20488 11796 20516
rect 11784 20479 11796 20488
rect 11790 20476 11796 20479
rect 11848 20476 11854 20528
rect 8122 20451 8180 20457
rect 8122 20448 8134 20451
rect 7800 20420 8134 20448
rect 7800 20408 7806 20420
rect 8122 20417 8134 20420
rect 8168 20417 8180 20451
rect 8122 20411 8180 20417
rect 8481 20451 8539 20457
rect 8481 20417 8493 20451
rect 8527 20417 8539 20451
rect 8481 20411 8539 20417
rect 8570 20408 8576 20460
rect 8628 20408 8634 20460
rect 9582 20408 9588 20460
rect 9640 20448 9646 20460
rect 13004 20457 13032 20556
rect 14458 20544 14464 20556
rect 14516 20544 14522 20596
rect 15841 20587 15899 20593
rect 15841 20553 15853 20587
rect 15887 20584 15899 20587
rect 17218 20584 17224 20596
rect 15887 20556 17224 20584
rect 15887 20553 15899 20556
rect 15841 20547 15899 20553
rect 17218 20544 17224 20556
rect 17276 20544 17282 20596
rect 15286 20516 15292 20528
rect 14660 20488 15292 20516
rect 10209 20451 10267 20457
rect 10209 20448 10221 20451
rect 9640 20420 10221 20448
rect 9640 20408 9646 20420
rect 10209 20417 10221 20420
rect 10255 20417 10267 20451
rect 10209 20411 10267 20417
rect 12989 20451 13047 20457
rect 12989 20417 13001 20451
rect 13035 20417 13047 20451
rect 13245 20451 13303 20457
rect 13245 20448 13257 20451
rect 12989 20411 13047 20417
rect 13096 20420 13257 20448
rect 8389 20383 8447 20389
rect 8389 20349 8401 20383
rect 8435 20380 8447 20383
rect 8588 20380 8616 20408
rect 8435 20352 8616 20380
rect 8435 20349 8447 20352
rect 8389 20343 8447 20349
rect 9950 20340 9956 20392
rect 10008 20340 10014 20392
rect 11514 20340 11520 20392
rect 11572 20340 11578 20392
rect 13096 20380 13124 20420
rect 13245 20417 13257 20420
rect 13291 20417 13303 20451
rect 13245 20411 13303 20417
rect 14461 20451 14519 20457
rect 14461 20417 14473 20451
rect 14507 20448 14519 20451
rect 14660 20448 14688 20488
rect 15286 20476 15292 20488
rect 15344 20476 15350 20528
rect 17672 20519 17730 20525
rect 17672 20485 17684 20519
rect 17718 20516 17730 20519
rect 18138 20516 18144 20528
rect 17718 20488 18144 20516
rect 17718 20485 17730 20488
rect 17672 20479 17730 20485
rect 18138 20476 18144 20488
rect 18196 20476 18202 20528
rect 18782 20476 18788 20528
rect 18840 20516 18846 20528
rect 19122 20519 19180 20525
rect 19122 20516 19134 20519
rect 18840 20488 19134 20516
rect 18840 20476 18846 20488
rect 19122 20485 19134 20488
rect 19168 20485 19180 20519
rect 19122 20479 19180 20485
rect 14507 20420 14688 20448
rect 14728 20451 14786 20457
rect 14507 20417 14519 20420
rect 14461 20411 14519 20417
rect 14728 20417 14740 20451
rect 14774 20448 14786 20451
rect 15194 20448 15200 20460
rect 14774 20420 15200 20448
rect 14774 20417 14786 20420
rect 14728 20411 14786 20417
rect 15194 20408 15200 20420
rect 15252 20408 15258 20460
rect 18046 20408 18052 20460
rect 18104 20448 18110 20460
rect 18877 20451 18935 20457
rect 18877 20448 18889 20451
rect 18104 20420 18889 20448
rect 18104 20408 18110 20420
rect 18877 20417 18889 20420
rect 18923 20417 18935 20451
rect 18877 20411 18935 20417
rect 12912 20352 13124 20380
rect 16025 20383 16083 20389
rect 6270 20272 6276 20324
rect 6328 20272 6334 20324
rect 12912 20321 12940 20352
rect 16025 20349 16037 20383
rect 16071 20349 16083 20383
rect 16025 20343 16083 20349
rect 12897 20315 12955 20321
rect 12897 20281 12909 20315
rect 12943 20281 12955 20315
rect 12897 20275 12955 20281
rect 14369 20315 14427 20321
rect 14369 20281 14381 20315
rect 14415 20312 14427 20315
rect 14458 20312 14464 20324
rect 14415 20284 14464 20312
rect 14415 20281 14427 20284
rect 14369 20275 14427 20281
rect 14458 20272 14464 20284
rect 14516 20272 14522 20324
rect 6181 20247 6239 20253
rect 6181 20213 6193 20247
rect 6227 20244 6239 20247
rect 6362 20244 6368 20256
rect 6227 20216 6368 20244
rect 6227 20213 6239 20216
rect 6181 20207 6239 20213
rect 6362 20204 6368 20216
rect 6420 20204 6426 20256
rect 6546 20204 6552 20256
rect 6604 20204 6610 20256
rect 7009 20247 7067 20253
rect 7009 20213 7021 20247
rect 7055 20244 7067 20247
rect 7650 20244 7656 20256
rect 7055 20216 7656 20244
rect 7055 20213 7067 20216
rect 7009 20207 7067 20213
rect 7650 20204 7656 20216
rect 7708 20204 7714 20256
rect 15102 20204 15108 20256
rect 15160 20244 15166 20256
rect 16040 20244 16068 20343
rect 16666 20340 16672 20392
rect 16724 20340 16730 20392
rect 17218 20340 17224 20392
rect 17276 20340 17282 20392
rect 17402 20340 17408 20392
rect 17460 20340 17466 20392
rect 16393 20315 16451 20321
rect 16393 20281 16405 20315
rect 16439 20312 16451 20315
rect 16684 20312 16712 20340
rect 16439 20284 16712 20312
rect 16439 20281 16451 20284
rect 16393 20275 16451 20281
rect 15160 20216 16068 20244
rect 15160 20204 15166 20216
rect 16482 20204 16488 20256
rect 16540 20204 16546 20256
rect 16666 20204 16672 20256
rect 16724 20204 16730 20256
rect 18785 20247 18843 20253
rect 18785 20213 18797 20247
rect 18831 20244 18843 20247
rect 19794 20244 19800 20256
rect 18831 20216 19800 20244
rect 18831 20213 18843 20216
rect 18785 20207 18843 20213
rect 19794 20204 19800 20216
rect 19852 20204 19858 20256
rect 20257 20247 20315 20253
rect 20257 20213 20269 20247
rect 20303 20244 20315 20247
rect 21450 20244 21456 20256
rect 20303 20216 21456 20244
rect 20303 20213 20315 20216
rect 20257 20207 20315 20213
rect 21450 20204 21456 20216
rect 21508 20204 21514 20256
rect 1104 20154 23828 20176
rect 1104 20102 1918 20154
rect 1970 20102 1982 20154
rect 2034 20102 2046 20154
rect 2098 20102 2110 20154
rect 2162 20102 2174 20154
rect 2226 20102 2238 20154
rect 2290 20102 7918 20154
rect 7970 20102 7982 20154
rect 8034 20102 8046 20154
rect 8098 20102 8110 20154
rect 8162 20102 8174 20154
rect 8226 20102 8238 20154
rect 8290 20102 13918 20154
rect 13970 20102 13982 20154
rect 14034 20102 14046 20154
rect 14098 20102 14110 20154
rect 14162 20102 14174 20154
rect 14226 20102 14238 20154
rect 14290 20102 19918 20154
rect 19970 20102 19982 20154
rect 20034 20102 20046 20154
rect 20098 20102 20110 20154
rect 20162 20102 20174 20154
rect 20226 20102 20238 20154
rect 20290 20102 23828 20154
rect 1104 20080 23828 20102
rect 5353 20043 5411 20049
rect 5353 20009 5365 20043
rect 5399 20040 5411 20043
rect 5626 20040 5632 20052
rect 5399 20012 5632 20040
rect 5399 20009 5411 20012
rect 5353 20003 5411 20009
rect 4709 19907 4767 19913
rect 4709 19873 4721 19907
rect 4755 19904 4767 19907
rect 5368 19904 5396 20003
rect 5626 20000 5632 20012
rect 5684 20000 5690 20052
rect 6546 20000 6552 20052
rect 6604 20040 6610 20052
rect 7009 20043 7067 20049
rect 6604 20012 6776 20040
rect 6604 20000 6610 20012
rect 6748 19913 6776 20012
rect 7009 20009 7021 20043
rect 7055 20040 7067 20043
rect 12437 20043 12495 20049
rect 7055 20012 9260 20040
rect 7055 20009 7067 20012
rect 7009 20003 7067 20009
rect 4755 19876 5396 19904
rect 6733 19907 6791 19913
rect 4755 19873 4767 19876
rect 4709 19867 4767 19873
rect 6733 19873 6745 19907
rect 6779 19873 6791 19907
rect 6733 19867 6791 19873
rect 8389 19907 8447 19913
rect 8389 19873 8401 19907
rect 8435 19904 8447 19907
rect 9122 19904 9128 19916
rect 8435 19876 9128 19904
rect 8435 19873 8447 19876
rect 8389 19867 8447 19873
rect 9122 19864 9128 19876
rect 9180 19864 9186 19916
rect 9232 19904 9260 20012
rect 9416 20012 12112 20040
rect 9416 19981 9444 20012
rect 9401 19975 9459 19981
rect 9401 19941 9413 19975
rect 9447 19941 9459 19975
rect 9401 19935 9459 19941
rect 9490 19932 9496 19984
rect 9548 19932 9554 19984
rect 9582 19932 9588 19984
rect 9640 19932 9646 19984
rect 9508 19904 9536 19932
rect 9232 19876 9536 19904
rect 10965 19907 11023 19913
rect 10965 19873 10977 19907
rect 11011 19904 11023 19907
rect 11011 19876 11192 19904
rect 11011 19873 11023 19876
rect 10965 19867 11023 19873
rect 8478 19836 8484 19848
rect 6288 19808 8484 19836
rect 6288 19780 6316 19808
rect 8478 19796 8484 19808
rect 8536 19796 8542 19848
rect 8570 19796 8576 19848
rect 8628 19796 8634 19848
rect 8662 19796 8668 19848
rect 8720 19836 8726 19848
rect 9033 19839 9091 19845
rect 9033 19836 9045 19839
rect 8720 19808 9045 19836
rect 8720 19796 8726 19808
rect 9033 19805 9045 19808
rect 9079 19836 9091 19839
rect 9306 19836 9312 19848
rect 9079 19808 9312 19836
rect 9079 19805 9091 19808
rect 9033 19799 9091 19805
rect 9306 19796 9312 19808
rect 9364 19796 9370 19848
rect 9490 19796 9496 19848
rect 9548 19796 9554 19848
rect 9858 19796 9864 19848
rect 9916 19836 9922 19848
rect 11057 19839 11115 19845
rect 11057 19836 11069 19839
rect 9916 19808 11069 19836
rect 9916 19796 9922 19808
rect 11057 19805 11069 19808
rect 11103 19805 11115 19839
rect 11164 19836 11192 19876
rect 11606 19836 11612 19848
rect 11164 19808 11612 19836
rect 11057 19799 11115 19805
rect 11606 19796 11612 19808
rect 11664 19796 11670 19848
rect 12084 19836 12112 20012
rect 12437 20009 12449 20043
rect 12483 20040 12495 20043
rect 12618 20040 12624 20052
rect 12483 20012 12624 20040
rect 12483 20009 12495 20012
rect 12437 20003 12495 20009
rect 12618 20000 12624 20012
rect 12676 20000 12682 20052
rect 12986 20000 12992 20052
rect 13044 20000 13050 20052
rect 14366 20000 14372 20052
rect 14424 20040 14430 20052
rect 15749 20043 15807 20049
rect 15749 20040 15761 20043
rect 14424 20012 15761 20040
rect 14424 20000 14430 20012
rect 15749 20009 15761 20012
rect 15795 20040 15807 20043
rect 17770 20040 17776 20052
rect 15795 20012 17776 20040
rect 15795 20009 15807 20012
rect 15749 20003 15807 20009
rect 17770 20000 17776 20012
rect 17828 20000 17834 20052
rect 12529 19975 12587 19981
rect 12529 19941 12541 19975
rect 12575 19972 12587 19975
rect 13004 19972 13032 20000
rect 12575 19944 13032 19972
rect 14461 19975 14519 19981
rect 12575 19941 12587 19944
rect 12529 19935 12587 19941
rect 14461 19941 14473 19975
rect 14507 19972 14519 19975
rect 15286 19972 15292 19984
rect 14507 19944 15292 19972
rect 14507 19941 14519 19944
rect 14461 19935 14519 19941
rect 15286 19932 15292 19944
rect 15344 19932 15350 19984
rect 12526 19836 12532 19848
rect 12084 19808 12532 19836
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 13262 19796 13268 19848
rect 13320 19836 13326 19848
rect 13642 19839 13700 19845
rect 13642 19836 13654 19839
rect 13320 19808 13654 19836
rect 13320 19796 13326 19808
rect 13642 19805 13654 19808
rect 13688 19805 13700 19839
rect 13642 19799 13700 19805
rect 13814 19796 13820 19848
rect 13872 19836 13878 19848
rect 13909 19839 13967 19845
rect 13909 19836 13921 19839
rect 13872 19808 13921 19836
rect 13872 19796 13878 19808
rect 13909 19805 13921 19808
rect 13955 19805 13967 19839
rect 13909 19799 13967 19805
rect 14277 19839 14335 19845
rect 14277 19805 14289 19839
rect 14323 19805 14335 19839
rect 14277 19799 14335 19805
rect 6270 19728 6276 19780
rect 6328 19728 6334 19780
rect 6362 19728 6368 19780
rect 6420 19768 6426 19780
rect 6466 19771 6524 19777
rect 6466 19768 6478 19771
rect 6420 19740 6478 19768
rect 6420 19728 6426 19740
rect 6466 19737 6478 19740
rect 6512 19737 6524 19771
rect 6466 19731 6524 19737
rect 7834 19728 7840 19780
rect 7892 19768 7898 19780
rect 8122 19771 8180 19777
rect 8122 19768 8134 19771
rect 7892 19740 8134 19768
rect 7892 19728 7898 19740
rect 8122 19737 8134 19740
rect 8168 19737 8180 19771
rect 8122 19731 8180 19737
rect 8294 19728 8300 19780
rect 8352 19768 8358 19780
rect 8588 19768 8616 19796
rect 8352 19740 8616 19768
rect 9125 19771 9183 19777
rect 8352 19728 8358 19740
rect 9125 19737 9137 19771
rect 9171 19737 9183 19771
rect 9125 19731 9183 19737
rect 10720 19771 10778 19777
rect 10720 19737 10732 19771
rect 10766 19768 10778 19771
rect 10870 19768 10876 19780
rect 10766 19740 10876 19768
rect 10766 19737 10778 19740
rect 10720 19731 10778 19737
rect 5258 19660 5264 19712
rect 5316 19660 5322 19712
rect 8570 19660 8576 19712
rect 8628 19660 8634 19712
rect 9140 19700 9168 19731
rect 10870 19728 10876 19740
rect 10928 19728 10934 19780
rect 11324 19771 11382 19777
rect 11324 19737 11336 19771
rect 11370 19768 11382 19771
rect 12066 19768 12072 19780
rect 11370 19740 12072 19768
rect 11370 19737 11382 19740
rect 11324 19731 11382 19737
rect 12066 19728 12072 19740
rect 12124 19728 12130 19780
rect 9674 19700 9680 19712
rect 9140 19672 9680 19700
rect 9674 19660 9680 19672
rect 9732 19660 9738 19712
rect 14292 19700 14320 19799
rect 14458 19796 14464 19848
rect 14516 19836 14522 19848
rect 14553 19839 14611 19845
rect 14553 19836 14565 19839
rect 14516 19808 14565 19836
rect 14516 19796 14522 19808
rect 14553 19805 14565 19808
rect 14599 19805 14611 19839
rect 14553 19799 14611 19805
rect 15194 19796 15200 19848
rect 15252 19796 15258 19848
rect 15470 19796 15476 19848
rect 15528 19836 15534 19848
rect 15528 19808 18460 19836
rect 15528 19796 15534 19808
rect 17034 19728 17040 19780
rect 17092 19728 17098 19780
rect 18046 19728 18052 19780
rect 18104 19768 18110 19780
rect 18242 19771 18300 19777
rect 18242 19768 18254 19771
rect 18104 19740 18254 19768
rect 18104 19728 18110 19740
rect 18242 19737 18254 19740
rect 18288 19737 18300 19771
rect 18432 19768 18460 19808
rect 18506 19796 18512 19848
rect 18564 19796 18570 19848
rect 18601 19839 18659 19845
rect 18601 19805 18613 19839
rect 18647 19805 18659 19839
rect 18601 19799 18659 19805
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19805 18935 19839
rect 18877 19799 18935 19805
rect 19245 19839 19303 19845
rect 19245 19805 19257 19839
rect 19291 19836 19303 19839
rect 19334 19836 19340 19848
rect 19291 19808 19340 19836
rect 19291 19805 19303 19808
rect 19245 19799 19303 19805
rect 18616 19768 18644 19799
rect 18432 19740 18644 19768
rect 18892 19768 18920 19799
rect 19334 19796 19340 19808
rect 19392 19796 19398 19848
rect 19518 19845 19524 19848
rect 19512 19836 19524 19845
rect 19479 19808 19524 19836
rect 19512 19799 19524 19808
rect 19518 19796 19524 19799
rect 19576 19796 19582 19848
rect 18892 19740 19380 19768
rect 18242 19731 18300 19737
rect 19352 19712 19380 19740
rect 14550 19700 14556 19712
rect 14292 19672 14556 19700
rect 14550 19660 14556 19672
rect 14608 19660 14614 19712
rect 17129 19703 17187 19709
rect 17129 19669 17141 19703
rect 17175 19700 17187 19703
rect 18138 19700 18144 19712
rect 17175 19672 18144 19700
rect 17175 19669 17187 19672
rect 17129 19663 17187 19669
rect 18138 19660 18144 19672
rect 18196 19660 18202 19712
rect 18690 19660 18696 19712
rect 18748 19660 18754 19712
rect 18966 19660 18972 19712
rect 19024 19660 19030 19712
rect 19334 19660 19340 19712
rect 19392 19660 19398 19712
rect 20625 19703 20683 19709
rect 20625 19669 20637 19703
rect 20671 19700 20683 19703
rect 21358 19700 21364 19712
rect 20671 19672 21364 19700
rect 20671 19669 20683 19672
rect 20625 19663 20683 19669
rect 21358 19660 21364 19672
rect 21416 19660 21422 19712
rect 1104 19610 23828 19632
rect 1104 19558 2658 19610
rect 2710 19558 2722 19610
rect 2774 19558 2786 19610
rect 2838 19558 2850 19610
rect 2902 19558 2914 19610
rect 2966 19558 2978 19610
rect 3030 19558 8658 19610
rect 8710 19558 8722 19610
rect 8774 19558 8786 19610
rect 8838 19558 8850 19610
rect 8902 19558 8914 19610
rect 8966 19558 8978 19610
rect 9030 19558 14658 19610
rect 14710 19558 14722 19610
rect 14774 19558 14786 19610
rect 14838 19558 14850 19610
rect 14902 19558 14914 19610
rect 14966 19558 14978 19610
rect 15030 19558 20658 19610
rect 20710 19558 20722 19610
rect 20774 19558 20786 19610
rect 20838 19558 20850 19610
rect 20902 19558 20914 19610
rect 20966 19558 20978 19610
rect 21030 19558 23828 19610
rect 1104 19536 23828 19558
rect 5258 19456 5264 19508
rect 5316 19496 5322 19508
rect 5316 19468 7144 19496
rect 5316 19456 5322 19468
rect 7006 19428 7012 19440
rect 6380 19400 7012 19428
rect 4614 19320 4620 19372
rect 4672 19360 4678 19372
rect 4709 19363 4767 19369
rect 4709 19360 4721 19363
rect 4672 19332 4721 19360
rect 4672 19320 4678 19332
rect 4709 19329 4721 19332
rect 4755 19329 4767 19363
rect 4709 19323 4767 19329
rect 4798 19320 4804 19372
rect 4856 19320 4862 19372
rect 5074 19369 5080 19372
rect 5068 19323 5080 19369
rect 5074 19320 5080 19323
rect 5132 19320 5138 19372
rect 6380 19369 6408 19400
rect 7006 19388 7012 19400
rect 7064 19388 7070 19440
rect 6365 19363 6423 19369
rect 6365 19329 6377 19363
rect 6411 19329 6423 19363
rect 6365 19323 6423 19329
rect 6457 19363 6515 19369
rect 6457 19329 6469 19363
rect 6503 19360 6515 19363
rect 6641 19363 6699 19369
rect 6641 19360 6653 19363
rect 6503 19332 6653 19360
rect 6503 19329 6515 19332
rect 6457 19323 6515 19329
rect 6641 19329 6653 19332
rect 6687 19329 6699 19363
rect 6641 19323 6699 19329
rect 6908 19363 6966 19369
rect 6908 19329 6920 19363
rect 6954 19360 6966 19363
rect 7116 19360 7144 19468
rect 7558 19456 7564 19508
rect 7616 19496 7622 19508
rect 8021 19499 8079 19505
rect 8021 19496 8033 19499
rect 7616 19468 8033 19496
rect 7616 19456 7622 19468
rect 8021 19465 8033 19468
rect 8067 19465 8079 19499
rect 8021 19459 8079 19465
rect 8386 19456 8392 19508
rect 8444 19456 8450 19508
rect 9490 19456 9496 19508
rect 9548 19496 9554 19508
rect 13722 19496 13728 19508
rect 9548 19468 13728 19496
rect 9548 19456 9554 19468
rect 13722 19456 13728 19468
rect 13780 19496 13786 19508
rect 14366 19496 14372 19508
rect 13780 19468 14372 19496
rect 13780 19456 13786 19468
rect 14366 19456 14372 19468
rect 14424 19456 14430 19508
rect 15194 19456 15200 19508
rect 15252 19496 15258 19508
rect 16485 19499 16543 19505
rect 16485 19496 16497 19499
rect 15252 19468 16497 19496
rect 15252 19456 15258 19468
rect 16485 19465 16497 19468
rect 16531 19465 16543 19499
rect 19797 19499 19855 19505
rect 19797 19496 19809 19499
rect 16485 19459 16543 19465
rect 16684 19468 19809 19496
rect 8404 19428 8432 19456
rect 12069 19431 12127 19437
rect 12069 19428 12081 19431
rect 8128 19400 8432 19428
rect 11624 19400 12081 19428
rect 8128 19369 8156 19400
rect 8386 19369 8392 19372
rect 6954 19332 7144 19360
rect 8113 19363 8171 19369
rect 6954 19329 6966 19332
rect 6908 19323 6966 19329
rect 8113 19329 8125 19363
rect 8159 19329 8171 19363
rect 8380 19360 8392 19369
rect 8347 19332 8392 19360
rect 8113 19323 8171 19329
rect 8380 19323 8392 19332
rect 8386 19320 8392 19323
rect 8444 19320 8450 19372
rect 9214 19320 9220 19372
rect 9272 19360 9278 19372
rect 9585 19363 9643 19369
rect 9585 19360 9597 19363
rect 9272 19332 9597 19360
rect 9272 19320 9278 19332
rect 9585 19329 9597 19332
rect 9631 19329 9643 19363
rect 9585 19323 9643 19329
rect 9852 19363 9910 19369
rect 9852 19329 9864 19363
rect 9898 19360 9910 19363
rect 10134 19360 10140 19372
rect 9898 19332 10140 19360
rect 9898 19329 9910 19332
rect 9852 19323 9910 19329
rect 10134 19320 10140 19332
rect 10192 19320 10198 19372
rect 10686 19320 10692 19372
rect 10744 19360 10750 19372
rect 11624 19369 11652 19400
rect 12069 19397 12081 19400
rect 12115 19397 12127 19431
rect 14461 19431 14519 19437
rect 14461 19428 14473 19431
rect 12069 19391 12127 19397
rect 12406 19400 14473 19428
rect 11333 19363 11391 19369
rect 11333 19360 11345 19363
rect 10744 19332 11345 19360
rect 10744 19320 10750 19332
rect 11333 19329 11345 19332
rect 11379 19329 11391 19363
rect 11333 19323 11391 19329
rect 11609 19363 11667 19369
rect 11609 19329 11621 19363
rect 11655 19329 11667 19363
rect 11609 19323 11667 19329
rect 10778 19252 10784 19304
rect 10836 19292 10842 19304
rect 10836 19264 11008 19292
rect 10836 19252 10842 19264
rect 10980 19233 11008 19264
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 11624 19292 11652 19323
rect 11698 19320 11704 19372
rect 11756 19320 11762 19372
rect 11112 19264 11652 19292
rect 11112 19252 11118 19264
rect 11882 19252 11888 19304
rect 11940 19292 11946 19304
rect 12406 19292 12434 19400
rect 14461 19397 14473 19400
rect 14507 19397 14519 19431
rect 14461 19391 14519 19397
rect 14820 19431 14878 19437
rect 14820 19397 14832 19431
rect 14866 19428 14878 19431
rect 16684 19428 16712 19468
rect 19797 19465 19809 19468
rect 19843 19465 19855 19499
rect 19797 19459 19855 19465
rect 21358 19456 21364 19508
rect 21416 19496 21422 19508
rect 21416 19468 22094 19496
rect 21416 19456 21422 19468
rect 14866 19400 16712 19428
rect 14866 19397 14878 19400
rect 14820 19391 14878 19397
rect 13170 19320 13176 19372
rect 13228 19360 13234 19372
rect 13817 19363 13875 19369
rect 13228 19332 13768 19360
rect 13228 19320 13234 19332
rect 11940 19264 12434 19292
rect 13740 19292 13768 19332
rect 13817 19329 13829 19363
rect 13863 19360 13875 19363
rect 14366 19360 14372 19372
rect 13863 19332 14372 19360
rect 13863 19329 13875 19332
rect 13817 19323 13875 19329
rect 14366 19320 14372 19332
rect 14424 19320 14430 19372
rect 14476 19360 14504 19391
rect 16758 19388 16764 19440
rect 16816 19428 16822 19440
rect 17402 19428 17408 19440
rect 16816 19400 17408 19428
rect 16816 19388 16822 19400
rect 17402 19388 17408 19400
rect 17460 19428 17466 19440
rect 19518 19428 19524 19440
rect 17460 19400 19524 19428
rect 17460 19388 17466 19400
rect 15102 19360 15108 19372
rect 14476 19332 15108 19360
rect 15102 19320 15108 19332
rect 15160 19360 15166 19372
rect 17218 19360 17224 19372
rect 15160 19332 15884 19360
rect 15160 19320 15166 19332
rect 14001 19295 14059 19301
rect 14001 19292 14013 19295
rect 13740 19264 14013 19292
rect 11940 19252 11946 19264
rect 14001 19261 14013 19264
rect 14047 19261 14059 19295
rect 14001 19255 14059 19261
rect 14550 19252 14556 19304
rect 14608 19252 14614 19304
rect 15856 19292 15884 19332
rect 16132 19332 17224 19360
rect 16025 19295 16083 19301
rect 16025 19292 16037 19295
rect 15856 19264 16037 19292
rect 16025 19261 16037 19264
rect 16071 19261 16083 19295
rect 16025 19255 16083 19261
rect 10965 19227 11023 19233
rect 10965 19193 10977 19227
rect 11011 19193 11023 19227
rect 10965 19187 11023 19193
rect 14185 19227 14243 19233
rect 14185 19193 14197 19227
rect 14231 19193 14243 19227
rect 14185 19187 14243 19193
rect 15933 19227 15991 19233
rect 15933 19193 15945 19227
rect 15979 19224 15991 19227
rect 16132 19224 16160 19332
rect 17218 19320 17224 19332
rect 17276 19320 17282 19372
rect 17977 19363 18035 19369
rect 17977 19329 17989 19363
rect 18023 19360 18035 19363
rect 18138 19360 18144 19372
rect 18023 19332 18144 19360
rect 18023 19329 18035 19332
rect 17977 19323 18035 19329
rect 18138 19320 18144 19332
rect 18196 19320 18202 19372
rect 18340 19369 18368 19400
rect 19518 19388 19524 19400
rect 19576 19388 19582 19440
rect 18325 19363 18383 19369
rect 18325 19329 18337 19363
rect 18371 19329 18383 19363
rect 18325 19323 18383 19329
rect 18414 19320 18420 19372
rect 18472 19360 18478 19372
rect 18581 19363 18639 19369
rect 18581 19360 18593 19363
rect 18472 19332 18593 19360
rect 18472 19320 18478 19332
rect 18581 19329 18593 19332
rect 18627 19329 18639 19363
rect 18581 19323 18639 19329
rect 19334 19320 19340 19372
rect 19392 19360 19398 19372
rect 20533 19363 20591 19369
rect 20533 19360 20545 19363
rect 19392 19332 20545 19360
rect 19392 19320 19398 19332
rect 20533 19329 20545 19332
rect 20579 19329 20591 19363
rect 22066 19360 22094 19468
rect 23017 19363 23075 19369
rect 23017 19360 23029 19363
rect 22066 19332 23029 19360
rect 20533 19323 20591 19329
rect 23017 19329 23029 19332
rect 23063 19329 23075 19363
rect 23017 19323 23075 19329
rect 23290 19320 23296 19372
rect 23348 19320 23354 19372
rect 18230 19252 18236 19304
rect 18288 19252 18294 19304
rect 18432 19292 18460 19320
rect 18340 19264 18460 19292
rect 15979 19196 16160 19224
rect 16393 19227 16451 19233
rect 15979 19193 15991 19196
rect 15933 19187 15991 19193
rect 16393 19193 16405 19227
rect 16439 19224 16451 19227
rect 16666 19224 16672 19236
rect 16439 19196 16672 19224
rect 16439 19193 16451 19196
rect 16393 19187 16451 19193
rect 4522 19116 4528 19168
rect 4580 19116 4586 19168
rect 5902 19116 5908 19168
rect 5960 19156 5966 19168
rect 6181 19159 6239 19165
rect 6181 19156 6193 19159
rect 5960 19128 6193 19156
rect 5960 19116 5966 19128
rect 6181 19125 6193 19128
rect 6227 19125 6239 19159
rect 6181 19119 6239 19125
rect 9493 19159 9551 19165
rect 9493 19125 9505 19159
rect 9539 19156 9551 19159
rect 9766 19156 9772 19168
rect 9539 19128 9772 19156
rect 9539 19125 9551 19128
rect 9493 19119 9551 19125
rect 9766 19116 9772 19128
rect 9824 19116 9830 19168
rect 10870 19116 10876 19168
rect 10928 19156 10934 19168
rect 11149 19159 11207 19165
rect 11149 19156 11161 19159
rect 10928 19128 11161 19156
rect 10928 19116 10934 19128
rect 11149 19125 11161 19128
rect 11195 19125 11207 19159
rect 14200 19156 14228 19187
rect 16666 19184 16672 19196
rect 16724 19184 16730 19236
rect 14918 19156 14924 19168
rect 14200 19128 14924 19156
rect 11149 19119 11207 19125
rect 14918 19116 14924 19128
rect 14976 19116 14982 19168
rect 16853 19159 16911 19165
rect 16853 19125 16865 19159
rect 16899 19156 16911 19159
rect 18340 19156 18368 19264
rect 20438 19252 20444 19304
rect 20496 19252 20502 19304
rect 19610 19184 19616 19236
rect 19668 19224 19674 19236
rect 20625 19227 20683 19233
rect 20625 19224 20637 19227
rect 19668 19196 20637 19224
rect 19668 19184 19674 19196
rect 20625 19193 20637 19196
rect 20671 19193 20683 19227
rect 20625 19187 20683 19193
rect 16899 19128 18368 19156
rect 16899 19125 16911 19128
rect 16853 19119 16911 19125
rect 19702 19116 19708 19168
rect 19760 19116 19766 19168
rect 1104 19066 23828 19088
rect 1104 19014 1918 19066
rect 1970 19014 1982 19066
rect 2034 19014 2046 19066
rect 2098 19014 2110 19066
rect 2162 19014 2174 19066
rect 2226 19014 2238 19066
rect 2290 19014 7918 19066
rect 7970 19014 7982 19066
rect 8034 19014 8046 19066
rect 8098 19014 8110 19066
rect 8162 19014 8174 19066
rect 8226 19014 8238 19066
rect 8290 19014 13918 19066
rect 13970 19014 13982 19066
rect 14034 19014 14046 19066
rect 14098 19014 14110 19066
rect 14162 19014 14174 19066
rect 14226 19014 14238 19066
rect 14290 19014 19918 19066
rect 19970 19014 19982 19066
rect 20034 19014 20046 19066
rect 20098 19014 20110 19066
rect 20162 19014 20174 19066
rect 20226 19014 20238 19066
rect 20290 19014 23828 19066
rect 1104 18992 23828 19014
rect 5074 18912 5080 18964
rect 5132 18952 5138 18964
rect 5261 18955 5319 18961
rect 5261 18952 5273 18955
rect 5132 18924 5273 18952
rect 5132 18912 5138 18924
rect 5261 18921 5273 18924
rect 5307 18921 5319 18955
rect 5261 18915 5319 18921
rect 6730 18912 6736 18964
rect 6788 18912 6794 18964
rect 8665 18955 8723 18961
rect 8665 18921 8677 18955
rect 8711 18952 8723 18955
rect 9858 18952 9864 18964
rect 8711 18924 9864 18952
rect 8711 18921 8723 18924
rect 8665 18915 8723 18921
rect 9858 18912 9864 18924
rect 9916 18912 9922 18964
rect 10042 18912 10048 18964
rect 10100 18912 10106 18964
rect 14185 18955 14243 18961
rect 14185 18921 14197 18955
rect 14231 18952 14243 18955
rect 14550 18952 14556 18964
rect 14231 18924 14556 18952
rect 14231 18921 14243 18924
rect 14185 18915 14243 18921
rect 14550 18912 14556 18924
rect 14608 18912 14614 18964
rect 18230 18912 18236 18964
rect 18288 18952 18294 18964
rect 18785 18955 18843 18961
rect 18785 18952 18797 18955
rect 18288 18924 18797 18952
rect 18288 18912 18294 18924
rect 18785 18921 18797 18924
rect 18831 18921 18843 18955
rect 18785 18915 18843 18921
rect 20438 18912 20444 18964
rect 20496 18952 20502 18964
rect 20625 18955 20683 18961
rect 20625 18952 20637 18955
rect 20496 18924 20637 18952
rect 20496 18912 20502 18924
rect 20625 18921 20637 18924
rect 20671 18921 20683 18955
rect 20625 18915 20683 18921
rect 8205 18887 8263 18893
rect 8205 18853 8217 18887
rect 8251 18884 8263 18887
rect 9582 18884 9588 18896
rect 8251 18856 9588 18884
rect 8251 18853 8263 18856
rect 8205 18847 8263 18853
rect 9582 18844 9588 18856
rect 9640 18844 9646 18896
rect 6822 18776 6828 18828
rect 6880 18776 6886 18828
rect 10060 18816 10088 18912
rect 15470 18884 15476 18896
rect 14568 18856 15476 18884
rect 7852 18788 10088 18816
rect 3878 18708 3884 18760
rect 3936 18708 3942 18760
rect 4148 18751 4206 18757
rect 4148 18717 4160 18751
rect 4194 18748 4206 18751
rect 4522 18748 4528 18760
rect 4194 18720 4528 18748
rect 4194 18717 4206 18720
rect 4148 18711 4206 18717
rect 4522 18708 4528 18720
rect 4580 18708 4586 18760
rect 5350 18708 5356 18760
rect 5408 18708 5414 18760
rect 5620 18751 5678 18757
rect 5620 18717 5632 18751
rect 5666 18748 5678 18751
rect 5902 18748 5908 18760
rect 5666 18720 5908 18748
rect 5666 18717 5678 18720
rect 5620 18711 5678 18717
rect 5902 18708 5908 18720
rect 5960 18708 5966 18760
rect 6914 18708 6920 18760
rect 6972 18748 6978 18760
rect 7081 18751 7139 18757
rect 7081 18748 7093 18751
rect 6972 18720 7093 18748
rect 6972 18708 6978 18720
rect 7081 18717 7093 18720
rect 7127 18717 7139 18751
rect 7081 18711 7139 18717
rect 4614 18640 4620 18692
rect 4672 18640 4678 18692
rect 5534 18640 5540 18692
rect 5592 18680 5598 18692
rect 7852 18680 7880 18788
rect 11514 18776 11520 18828
rect 11572 18816 11578 18828
rect 11793 18819 11851 18825
rect 11793 18816 11805 18819
rect 11572 18788 11805 18816
rect 11572 18776 11578 18788
rect 11793 18785 11805 18788
rect 11839 18785 11851 18819
rect 14568 18816 14596 18856
rect 15470 18844 15476 18856
rect 15528 18884 15534 18896
rect 15933 18887 15991 18893
rect 15933 18884 15945 18887
rect 15528 18856 15945 18884
rect 15528 18844 15534 18856
rect 15933 18853 15945 18856
rect 15979 18853 15991 18887
rect 15933 18847 15991 18853
rect 16485 18887 16543 18893
rect 16485 18853 16497 18887
rect 16531 18853 16543 18887
rect 16485 18847 16543 18853
rect 11793 18779 11851 18785
rect 14108 18788 14596 18816
rect 8478 18708 8484 18760
rect 8536 18748 8542 18760
rect 8573 18751 8631 18757
rect 8573 18748 8585 18751
rect 8536 18720 8585 18748
rect 8536 18708 8542 18720
rect 8573 18717 8585 18720
rect 8619 18748 8631 18751
rect 10502 18748 10508 18760
rect 8619 18720 10508 18748
rect 8619 18717 8631 18720
rect 8573 18711 8631 18717
rect 10502 18708 10508 18720
rect 10560 18708 10566 18760
rect 10962 18708 10968 18760
rect 11020 18708 11026 18760
rect 11146 18708 11152 18760
rect 11204 18708 11210 18760
rect 11808 18748 11836 18779
rect 11808 18720 12434 18748
rect 5592 18652 7880 18680
rect 8941 18683 8999 18689
rect 5592 18640 5598 18652
rect 8941 18649 8953 18683
rect 8987 18680 8999 18683
rect 9490 18680 9496 18692
rect 8987 18652 9496 18680
rect 8987 18649 8999 18652
rect 8941 18643 8999 18649
rect 9490 18640 9496 18652
rect 9548 18640 9554 18692
rect 12060 18683 12118 18689
rect 12060 18649 12072 18683
rect 12106 18649 12118 18683
rect 12406 18680 12434 18720
rect 13354 18708 13360 18760
rect 13412 18708 13418 18760
rect 14108 18757 14136 18788
rect 14568 18760 14596 18788
rect 14642 18776 14648 18828
rect 14700 18816 14706 18828
rect 15194 18816 15200 18828
rect 14700 18788 15200 18816
rect 14700 18776 14706 18788
rect 15194 18776 15200 18788
rect 15252 18776 15258 18828
rect 14093 18751 14151 18757
rect 14093 18717 14105 18751
rect 14139 18717 14151 18751
rect 14093 18711 14151 18717
rect 14369 18751 14427 18757
rect 14369 18717 14381 18751
rect 14415 18748 14427 18751
rect 14458 18748 14464 18760
rect 14415 18720 14464 18748
rect 14415 18717 14427 18720
rect 14369 18711 14427 18717
rect 14458 18708 14464 18720
rect 14516 18708 14522 18760
rect 14550 18708 14556 18760
rect 14608 18708 14614 18760
rect 16500 18748 16528 18847
rect 17865 18819 17923 18825
rect 17865 18785 17877 18819
rect 17911 18816 17923 18819
rect 18690 18816 18696 18828
rect 17911 18788 18696 18816
rect 17911 18785 17923 18788
rect 17865 18779 17923 18785
rect 18690 18776 18696 18788
rect 18748 18776 18754 18828
rect 18966 18776 18972 18828
rect 19024 18816 19030 18828
rect 19245 18819 19303 18825
rect 19245 18816 19257 18819
rect 19024 18788 19257 18816
rect 19024 18776 19030 18788
rect 19245 18785 19257 18788
rect 19291 18785 19303 18819
rect 19245 18779 19303 18785
rect 18509 18751 18567 18757
rect 18509 18748 18521 18751
rect 16500 18720 18521 18748
rect 18509 18717 18521 18720
rect 18555 18717 18567 18751
rect 18509 18711 18567 18717
rect 18874 18708 18880 18760
rect 18932 18708 18938 18760
rect 20717 18751 20775 18757
rect 20717 18748 20729 18751
rect 19168 18720 20729 18748
rect 13814 18680 13820 18692
rect 12406 18652 13820 18680
rect 12060 18643 12118 18649
rect 4632 18612 4660 18640
rect 10042 18612 10048 18624
rect 4632 18584 10048 18612
rect 10042 18572 10048 18584
rect 10100 18572 10106 18624
rect 10873 18615 10931 18621
rect 10873 18581 10885 18615
rect 10919 18612 10931 18615
rect 11422 18612 11428 18624
rect 10919 18584 11428 18612
rect 10919 18581 10931 18584
rect 10873 18575 10931 18581
rect 11422 18572 11428 18584
rect 11480 18572 11486 18624
rect 11701 18615 11759 18621
rect 11701 18581 11713 18615
rect 11747 18612 11759 18615
rect 11790 18612 11796 18624
rect 11747 18584 11796 18612
rect 11747 18581 11759 18584
rect 11701 18575 11759 18581
rect 11790 18572 11796 18584
rect 11848 18572 11854 18624
rect 11974 18572 11980 18624
rect 12032 18612 12038 18624
rect 12084 18612 12112 18643
rect 13814 18640 13820 18652
rect 13872 18640 13878 18692
rect 13998 18640 14004 18692
rect 14056 18680 14062 18692
rect 14645 18683 14703 18689
rect 14645 18680 14657 18683
rect 14056 18652 14657 18680
rect 14056 18640 14062 18652
rect 14645 18649 14657 18652
rect 14691 18649 14703 18683
rect 14645 18643 14703 18649
rect 17620 18683 17678 18689
rect 17620 18649 17632 18683
rect 17666 18680 17678 18683
rect 19168 18680 19196 18720
rect 20717 18717 20729 18720
rect 20763 18717 20775 18751
rect 20717 18711 20775 18717
rect 21266 18708 21272 18760
rect 21324 18708 21330 18760
rect 21450 18708 21456 18760
rect 21508 18748 21514 18760
rect 23017 18751 23075 18757
rect 23017 18748 23029 18751
rect 21508 18720 23029 18748
rect 21508 18708 21514 18720
rect 23017 18717 23029 18720
rect 23063 18717 23075 18751
rect 23017 18711 23075 18717
rect 17666 18652 19196 18680
rect 19512 18683 19570 18689
rect 17666 18649 17678 18652
rect 17620 18643 17678 18649
rect 19512 18649 19524 18683
rect 19558 18680 19570 18683
rect 19794 18680 19800 18692
rect 19558 18652 19800 18680
rect 19558 18649 19570 18652
rect 19512 18643 19570 18649
rect 19794 18640 19800 18652
rect 19852 18640 19858 18692
rect 23290 18640 23296 18692
rect 23348 18640 23354 18692
rect 12032 18584 12112 18612
rect 12032 18572 12038 18584
rect 13170 18572 13176 18624
rect 13228 18572 13234 18624
rect 13538 18572 13544 18624
rect 13596 18612 13602 18624
rect 13909 18615 13967 18621
rect 13909 18612 13921 18615
rect 13596 18584 13921 18612
rect 13596 18572 13602 18584
rect 13909 18581 13921 18584
rect 13955 18581 13967 18615
rect 13909 18575 13967 18581
rect 14274 18572 14280 18624
rect 14332 18612 14338 18624
rect 14553 18615 14611 18621
rect 14553 18612 14565 18615
rect 14332 18584 14565 18612
rect 14332 18572 14338 18584
rect 14553 18581 14565 18584
rect 14599 18581 14611 18615
rect 14553 18575 14611 18581
rect 17954 18572 17960 18624
rect 18012 18572 18018 18624
rect 1104 18522 23828 18544
rect 1104 18470 2658 18522
rect 2710 18470 2722 18522
rect 2774 18470 2786 18522
rect 2838 18470 2850 18522
rect 2902 18470 2914 18522
rect 2966 18470 2978 18522
rect 3030 18470 8658 18522
rect 8710 18470 8722 18522
rect 8774 18470 8786 18522
rect 8838 18470 8850 18522
rect 8902 18470 8914 18522
rect 8966 18470 8978 18522
rect 9030 18470 14658 18522
rect 14710 18470 14722 18522
rect 14774 18470 14786 18522
rect 14838 18470 14850 18522
rect 14902 18470 14914 18522
rect 14966 18470 14978 18522
rect 15030 18470 20658 18522
rect 20710 18470 20722 18522
rect 20774 18470 20786 18522
rect 20838 18470 20850 18522
rect 20902 18470 20914 18522
rect 20966 18470 20978 18522
rect 21030 18470 23828 18522
rect 1104 18448 23828 18470
rect 3878 18368 3884 18420
rect 3936 18408 3942 18420
rect 4065 18411 4123 18417
rect 4065 18408 4077 18411
rect 3936 18380 4077 18408
rect 3936 18368 3942 18380
rect 4065 18377 4077 18380
rect 4111 18377 4123 18411
rect 4065 18371 4123 18377
rect 4341 18411 4399 18417
rect 4341 18377 4353 18411
rect 4387 18408 4399 18411
rect 5350 18408 5356 18420
rect 4387 18380 5356 18408
rect 4387 18377 4399 18380
rect 4341 18371 4399 18377
rect 5350 18368 5356 18380
rect 5408 18368 5414 18420
rect 5442 18368 5448 18420
rect 5500 18408 5506 18420
rect 5500 18380 6408 18408
rect 5500 18368 5506 18380
rect 6270 18340 6276 18352
rect 4448 18312 6276 18340
rect 4154 18232 4160 18284
rect 4212 18232 4218 18284
rect 4448 18281 4476 18312
rect 6270 18300 6276 18312
rect 6328 18300 6334 18352
rect 6380 18340 6408 18380
rect 9306 18368 9312 18420
rect 9364 18408 9370 18420
rect 9861 18411 9919 18417
rect 9861 18408 9873 18411
rect 9364 18380 9873 18408
rect 9364 18368 9370 18380
rect 9861 18377 9873 18380
rect 9907 18377 9919 18411
rect 9861 18371 9919 18377
rect 10042 18368 10048 18420
rect 10100 18408 10106 18420
rect 11517 18411 11575 18417
rect 11517 18408 11529 18411
rect 10100 18380 11529 18408
rect 10100 18368 10106 18380
rect 11517 18377 11529 18380
rect 11563 18377 11575 18411
rect 11517 18371 11575 18377
rect 13998 18368 14004 18420
rect 14056 18368 14062 18420
rect 14366 18368 14372 18420
rect 14424 18408 14430 18420
rect 15102 18408 15108 18420
rect 14424 18380 15108 18408
rect 14424 18368 14430 18380
rect 15102 18368 15108 18380
rect 15160 18408 15166 18420
rect 15289 18411 15347 18417
rect 15289 18408 15301 18411
rect 15160 18380 15301 18408
rect 15160 18368 15166 18380
rect 15289 18377 15301 18380
rect 15335 18377 15347 18411
rect 15289 18371 15347 18377
rect 18046 18368 18052 18420
rect 18104 18368 18110 18420
rect 18138 18368 18144 18420
rect 18196 18368 18202 18420
rect 20993 18411 21051 18417
rect 20993 18377 21005 18411
rect 21039 18408 21051 18411
rect 21266 18408 21272 18420
rect 21039 18380 21272 18408
rect 21039 18377 21051 18380
rect 20993 18371 21051 18377
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 6886 18343 6944 18349
rect 6886 18340 6898 18343
rect 6380 18312 6898 18340
rect 6886 18309 6898 18312
rect 6932 18309 6944 18343
rect 6886 18303 6944 18309
rect 11333 18343 11391 18349
rect 11333 18309 11345 18343
rect 11379 18340 11391 18343
rect 13909 18343 13967 18349
rect 13909 18340 13921 18343
rect 11379 18312 13921 18340
rect 11379 18309 11391 18312
rect 11333 18303 11391 18309
rect 13909 18309 13921 18312
rect 13955 18340 13967 18343
rect 14016 18340 14044 18368
rect 13955 18312 14044 18340
rect 13955 18309 13967 18312
rect 13909 18303 13967 18309
rect 16850 18300 16856 18352
rect 16908 18340 16914 18352
rect 19254 18343 19312 18349
rect 19254 18340 19266 18343
rect 16908 18312 19266 18340
rect 16908 18300 16914 18312
rect 19254 18309 19266 18312
rect 19300 18309 19312 18343
rect 19254 18303 19312 18309
rect 19702 18300 19708 18352
rect 19760 18340 19766 18352
rect 19858 18343 19916 18349
rect 19858 18340 19870 18343
rect 19760 18312 19870 18340
rect 19760 18300 19766 18312
rect 19858 18309 19870 18312
rect 19904 18309 19916 18343
rect 19858 18303 19916 18309
rect 4433 18275 4491 18281
rect 4433 18241 4445 18275
rect 4479 18241 4491 18275
rect 4433 18235 4491 18241
rect 4525 18275 4583 18281
rect 4525 18241 4537 18275
rect 4571 18272 4583 18275
rect 5534 18272 5540 18284
rect 4571 18244 5540 18272
rect 4571 18241 4583 18244
rect 4525 18235 4583 18241
rect 5534 18232 5540 18244
rect 5592 18232 5598 18284
rect 5925 18275 5983 18281
rect 5925 18241 5937 18275
rect 5971 18272 5983 18275
rect 6086 18272 6092 18284
rect 5971 18244 6092 18272
rect 5971 18241 5983 18244
rect 5925 18235 5983 18241
rect 6086 18232 6092 18244
rect 6144 18232 6150 18284
rect 6178 18232 6184 18284
rect 6236 18232 6242 18284
rect 6549 18275 6607 18281
rect 6549 18241 6561 18275
rect 6595 18272 6607 18275
rect 6730 18272 6736 18284
rect 6595 18244 6736 18272
rect 6595 18241 6607 18244
rect 6549 18235 6607 18241
rect 6730 18232 6736 18244
rect 6788 18232 6794 18284
rect 7466 18232 7472 18284
rect 7524 18272 7530 18284
rect 9226 18275 9284 18281
rect 9226 18272 9238 18275
rect 7524 18244 9238 18272
rect 7524 18232 7530 18244
rect 9226 18241 9238 18244
rect 9272 18241 9284 18275
rect 9226 18235 9284 18241
rect 10594 18232 10600 18284
rect 10652 18272 10658 18284
rect 12161 18275 12219 18281
rect 12161 18272 12173 18275
rect 10652 18244 12173 18272
rect 10652 18232 10658 18244
rect 12161 18241 12173 18244
rect 12207 18241 12219 18275
rect 12161 18235 12219 18241
rect 14001 18275 14059 18281
rect 14001 18241 14013 18275
rect 14047 18272 14059 18275
rect 14458 18272 14464 18284
rect 14047 18244 14464 18272
rect 14047 18241 14059 18244
rect 14001 18235 14059 18241
rect 14458 18232 14464 18244
rect 14516 18232 14522 18284
rect 16669 18275 16727 18281
rect 16669 18241 16681 18275
rect 16715 18272 16727 18275
rect 16758 18272 16764 18284
rect 16715 18244 16764 18272
rect 16715 18241 16727 18244
rect 16669 18235 16727 18241
rect 16758 18232 16764 18244
rect 16816 18232 16822 18284
rect 16942 18281 16948 18284
rect 16936 18235 16948 18281
rect 16942 18232 16948 18235
rect 17000 18232 17006 18284
rect 4890 18164 4896 18216
rect 4948 18164 4954 18216
rect 6196 18204 6224 18232
rect 6641 18207 6699 18213
rect 6641 18204 6653 18207
rect 6196 18176 6653 18204
rect 6641 18173 6653 18176
rect 6687 18173 6699 18207
rect 6641 18167 6699 18173
rect 9493 18207 9551 18213
rect 9493 18173 9505 18207
rect 9539 18204 9551 18207
rect 9858 18204 9864 18216
rect 9539 18176 9864 18204
rect 9539 18173 9551 18176
rect 9493 18167 9551 18173
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 11882 18164 11888 18216
rect 11940 18204 11946 18216
rect 11977 18207 12035 18213
rect 11977 18204 11989 18207
rect 11940 18176 11989 18204
rect 11940 18164 11946 18176
rect 11977 18173 11989 18176
rect 12023 18173 12035 18207
rect 11977 18167 12035 18173
rect 13262 18164 13268 18216
rect 13320 18204 13326 18216
rect 16393 18207 16451 18213
rect 16393 18204 16405 18207
rect 13320 18176 16405 18204
rect 13320 18164 13326 18176
rect 16393 18173 16405 18176
rect 16439 18173 16451 18207
rect 16393 18167 16451 18173
rect 19518 18164 19524 18216
rect 19576 18164 19582 18216
rect 19610 18164 19616 18216
rect 19668 18164 19674 18216
rect 4709 18139 4767 18145
rect 4709 18105 4721 18139
rect 4755 18136 4767 18139
rect 4908 18136 4936 18164
rect 4755 18108 4936 18136
rect 4755 18105 4767 18108
rect 4709 18099 4767 18105
rect 7834 18096 7840 18148
rect 7892 18136 7898 18148
rect 8113 18139 8171 18145
rect 8113 18136 8125 18139
rect 7892 18108 8125 18136
rect 7892 18096 7898 18108
rect 8113 18105 8125 18108
rect 8159 18105 8171 18139
rect 8113 18099 8171 18105
rect 11238 18096 11244 18148
rect 11296 18136 11302 18148
rect 11609 18139 11667 18145
rect 11609 18136 11621 18139
rect 11296 18108 11621 18136
rect 11296 18096 11302 18108
rect 11609 18105 11621 18108
rect 11655 18105 11667 18139
rect 11609 18099 11667 18105
rect 14642 18096 14648 18148
rect 14700 18136 14706 18148
rect 15194 18136 15200 18148
rect 14700 18108 15200 18136
rect 14700 18096 14706 18108
rect 15194 18096 15200 18108
rect 15252 18096 15258 18148
rect 4801 18071 4859 18077
rect 4801 18037 4813 18071
rect 4847 18068 4859 18071
rect 4890 18068 4896 18080
rect 4847 18040 4896 18068
rect 4847 18037 4859 18040
rect 4801 18031 4859 18037
rect 4890 18028 4896 18040
rect 4948 18028 4954 18080
rect 6270 18028 6276 18080
rect 6328 18068 6334 18080
rect 6365 18071 6423 18077
rect 6365 18068 6377 18071
rect 6328 18040 6377 18068
rect 6328 18028 6334 18040
rect 6365 18037 6377 18040
rect 6411 18037 6423 18071
rect 6365 18031 6423 18037
rect 8021 18071 8079 18077
rect 8021 18037 8033 18071
rect 8067 18068 8079 18071
rect 8386 18068 8392 18080
rect 8067 18040 8392 18068
rect 8067 18037 8079 18040
rect 8021 18031 8079 18037
rect 8386 18028 8392 18040
rect 8444 18028 8450 18080
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 15841 18071 15899 18077
rect 15841 18068 15853 18071
rect 14792 18040 15853 18068
rect 14792 18028 14798 18040
rect 15841 18037 15853 18040
rect 15887 18037 15899 18071
rect 15841 18031 15899 18037
rect 1104 17978 23828 18000
rect 1104 17926 1918 17978
rect 1970 17926 1982 17978
rect 2034 17926 2046 17978
rect 2098 17926 2110 17978
rect 2162 17926 2174 17978
rect 2226 17926 2238 17978
rect 2290 17926 7918 17978
rect 7970 17926 7982 17978
rect 8034 17926 8046 17978
rect 8098 17926 8110 17978
rect 8162 17926 8174 17978
rect 8226 17926 8238 17978
rect 8290 17926 13918 17978
rect 13970 17926 13982 17978
rect 14034 17926 14046 17978
rect 14098 17926 14110 17978
rect 14162 17926 14174 17978
rect 14226 17926 14238 17978
rect 14290 17926 19918 17978
rect 19970 17926 19982 17978
rect 20034 17926 20046 17978
rect 20098 17926 20110 17978
rect 20162 17926 20174 17978
rect 20226 17926 20238 17978
rect 20290 17926 23828 17978
rect 1104 17904 23828 17926
rect 7466 17864 7472 17876
rect 3896 17836 7472 17864
rect 3896 17660 3924 17836
rect 7466 17824 7472 17836
rect 7524 17824 7530 17876
rect 9125 17867 9183 17873
rect 9125 17833 9137 17867
rect 9171 17864 9183 17867
rect 10594 17864 10600 17876
rect 9171 17836 10600 17864
rect 9171 17833 9183 17836
rect 9125 17827 9183 17833
rect 10594 17824 10600 17836
rect 10652 17824 10658 17876
rect 11146 17824 11152 17876
rect 11204 17864 11210 17876
rect 11333 17867 11391 17873
rect 11333 17864 11345 17867
rect 11204 17836 11345 17864
rect 11204 17824 11210 17836
rect 11333 17833 11345 17836
rect 11379 17833 11391 17867
rect 11333 17827 11391 17833
rect 13354 17824 13360 17876
rect 13412 17864 13418 17876
rect 13449 17867 13507 17873
rect 13449 17864 13461 17867
rect 13412 17836 13461 17864
rect 13412 17824 13418 17836
rect 13449 17833 13461 17836
rect 13495 17833 13507 17867
rect 13449 17827 13507 17833
rect 14553 17867 14611 17873
rect 14553 17833 14565 17867
rect 14599 17864 14611 17867
rect 14642 17864 14648 17876
rect 14599 17836 14648 17864
rect 14599 17833 14611 17836
rect 14553 17827 14611 17833
rect 14642 17824 14648 17836
rect 14700 17824 14706 17876
rect 16117 17867 16175 17873
rect 14752 17836 15700 17864
rect 4706 17756 4712 17808
rect 4764 17796 4770 17808
rect 4764 17768 8892 17796
rect 4764 17756 4770 17768
rect 4246 17688 4252 17740
rect 4304 17728 4310 17740
rect 7006 17728 7012 17740
rect 4304 17700 7012 17728
rect 4304 17688 4310 17700
rect 7006 17688 7012 17700
rect 7064 17688 7070 17740
rect 4065 17663 4123 17669
rect 4065 17660 4077 17663
rect 3896 17632 4077 17660
rect 4065 17629 4077 17632
rect 4111 17629 4123 17663
rect 4065 17623 4123 17629
rect 4709 17663 4767 17669
rect 4709 17629 4721 17663
rect 4755 17660 4767 17663
rect 5350 17660 5356 17672
rect 4755 17632 5356 17660
rect 4755 17629 4767 17632
rect 4709 17623 4767 17629
rect 5350 17620 5356 17632
rect 5408 17620 5414 17672
rect 6917 17663 6975 17669
rect 6917 17629 6929 17663
rect 6963 17629 6975 17663
rect 6917 17623 6975 17629
rect 4801 17595 4859 17601
rect 4801 17561 4813 17595
rect 4847 17561 4859 17595
rect 4801 17555 4859 17561
rect 3510 17484 3516 17536
rect 3568 17524 3574 17536
rect 4154 17524 4160 17536
rect 3568 17496 4160 17524
rect 3568 17484 3574 17496
rect 4154 17484 4160 17496
rect 4212 17524 4218 17536
rect 4816 17524 4844 17555
rect 6546 17552 6552 17604
rect 6604 17552 6610 17604
rect 6932 17536 6960 17623
rect 8478 17552 8484 17604
rect 8536 17592 8542 17604
rect 8757 17595 8815 17601
rect 8757 17592 8769 17595
rect 8536 17564 8769 17592
rect 8536 17552 8542 17564
rect 8757 17561 8769 17564
rect 8803 17561 8815 17595
rect 8864 17592 8892 17768
rect 11606 17756 11612 17808
rect 11664 17756 11670 17808
rect 14461 17799 14519 17805
rect 14461 17765 14473 17799
rect 14507 17796 14519 17799
rect 14752 17796 14780 17836
rect 14507 17768 14780 17796
rect 15672 17796 15700 17836
rect 16117 17833 16129 17867
rect 16163 17864 16175 17867
rect 16942 17864 16948 17876
rect 16163 17836 16948 17864
rect 16163 17833 16175 17836
rect 16117 17827 16175 17833
rect 16942 17824 16948 17836
rect 17000 17824 17006 17876
rect 18506 17824 18512 17876
rect 18564 17864 18570 17876
rect 18693 17867 18751 17873
rect 18693 17864 18705 17867
rect 18564 17836 18705 17864
rect 18564 17824 18570 17836
rect 18693 17833 18705 17836
rect 18739 17833 18751 17867
rect 18693 17827 18751 17833
rect 17954 17796 17960 17808
rect 15672 17768 17960 17796
rect 14507 17765 14519 17768
rect 14461 17759 14519 17765
rect 17954 17756 17960 17768
rect 18012 17756 18018 17808
rect 18874 17756 18880 17808
rect 18932 17756 18938 17808
rect 9674 17688 9680 17740
rect 9732 17728 9738 17740
rect 9953 17731 10011 17737
rect 9953 17728 9965 17731
rect 9732 17700 9965 17728
rect 9732 17688 9738 17700
rect 9953 17697 9965 17700
rect 9999 17697 10011 17731
rect 9953 17691 10011 17697
rect 11517 17731 11575 17737
rect 11517 17697 11529 17731
rect 11563 17697 11575 17731
rect 11517 17691 11575 17697
rect 8941 17663 8999 17669
rect 8941 17629 8953 17663
rect 8987 17660 8999 17663
rect 9122 17660 9128 17672
rect 8987 17632 9128 17660
rect 8987 17629 8999 17632
rect 8941 17623 8999 17629
rect 9122 17620 9128 17632
rect 9180 17620 9186 17672
rect 9309 17663 9367 17669
rect 9309 17629 9321 17663
rect 9355 17660 9367 17663
rect 11532 17660 11560 17691
rect 11698 17688 11704 17740
rect 11756 17728 11762 17740
rect 12069 17731 12127 17737
rect 12069 17728 12081 17731
rect 11756 17700 12081 17728
rect 11756 17688 11762 17700
rect 12069 17697 12081 17700
rect 12115 17697 12127 17731
rect 18417 17731 18475 17737
rect 18417 17728 18429 17731
rect 12069 17691 12127 17697
rect 16592 17700 18429 17728
rect 9355 17632 11560 17660
rect 9355 17629 9367 17632
rect 9309 17623 9367 17629
rect 11882 17620 11888 17672
rect 11940 17660 11946 17672
rect 11977 17663 12035 17669
rect 11977 17660 11989 17663
rect 11940 17632 11989 17660
rect 11940 17620 11946 17632
rect 11977 17629 11989 17632
rect 12023 17660 12035 17663
rect 12023 17632 12434 17660
rect 12023 17629 12035 17632
rect 11977 17623 12035 17629
rect 10198 17595 10256 17601
rect 10198 17592 10210 17595
rect 8864 17564 10210 17592
rect 8757 17555 8815 17561
rect 10198 17561 10210 17564
rect 10244 17561 10256 17595
rect 10198 17555 10256 17561
rect 10686 17552 10692 17604
rect 10744 17552 10750 17604
rect 12066 17552 12072 17604
rect 12124 17592 12130 17604
rect 12314 17595 12372 17601
rect 12314 17592 12326 17595
rect 12124 17564 12326 17592
rect 12124 17552 12130 17564
rect 12314 17561 12326 17564
rect 12360 17561 12372 17595
rect 12406 17592 12434 17632
rect 13722 17620 13728 17672
rect 13780 17620 13786 17672
rect 14093 17663 14151 17669
rect 14093 17629 14105 17663
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 14108 17592 14136 17623
rect 14366 17620 14372 17672
rect 14424 17620 14430 17672
rect 14737 17663 14795 17669
rect 14737 17629 14749 17663
rect 14783 17660 14795 17663
rect 16592 17660 16620 17700
rect 18417 17697 18429 17700
rect 18463 17697 18475 17731
rect 18892 17728 18920 17756
rect 18417 17691 18475 17697
rect 18800 17700 18920 17728
rect 14783 17632 16620 17660
rect 14783 17629 14795 17632
rect 14737 17623 14795 17629
rect 18046 17620 18052 17672
rect 18104 17660 18110 17672
rect 18800 17669 18828 17700
rect 18233 17663 18291 17669
rect 18233 17660 18245 17663
rect 18104 17632 18245 17660
rect 18104 17620 18110 17632
rect 18233 17629 18245 17632
rect 18279 17660 18291 17663
rect 18509 17663 18567 17669
rect 18509 17660 18521 17663
rect 18279 17632 18521 17660
rect 18279 17629 18291 17632
rect 18233 17623 18291 17629
rect 18509 17629 18521 17632
rect 18555 17629 18567 17663
rect 18509 17623 18567 17629
rect 18785 17663 18843 17669
rect 18785 17629 18797 17663
rect 18831 17629 18843 17663
rect 18785 17623 18843 17629
rect 18877 17663 18935 17669
rect 18877 17629 18889 17663
rect 18923 17660 18935 17663
rect 19058 17660 19064 17672
rect 18923 17632 19064 17660
rect 18923 17629 18935 17632
rect 18877 17623 18935 17629
rect 19058 17620 19064 17632
rect 19116 17620 19122 17672
rect 19334 17620 19340 17672
rect 19392 17620 19398 17672
rect 12406 17564 14136 17592
rect 14384 17592 14412 17620
rect 14982 17595 15040 17601
rect 14982 17592 14994 17595
rect 14384 17564 14994 17592
rect 12314 17555 12372 17561
rect 14982 17561 14994 17564
rect 15028 17561 15040 17595
rect 14982 17555 15040 17561
rect 15102 17552 15108 17604
rect 15160 17592 15166 17604
rect 16209 17595 16267 17601
rect 16209 17592 16221 17595
rect 15160 17564 16221 17592
rect 15160 17552 15166 17564
rect 16209 17561 16221 17564
rect 16255 17561 16267 17595
rect 19352 17592 19380 17620
rect 16209 17555 16267 17561
rect 17512 17564 19380 17592
rect 4212 17496 4844 17524
rect 4212 17484 4218 17496
rect 6822 17484 6828 17536
rect 6880 17484 6886 17536
rect 6914 17484 6920 17536
rect 6972 17484 6978 17536
rect 9861 17527 9919 17533
rect 9861 17493 9873 17527
rect 9907 17524 9919 17527
rect 10704 17524 10732 17552
rect 9907 17496 10732 17524
rect 9907 17493 9919 17496
rect 9861 17487 9919 17493
rect 13630 17484 13636 17536
rect 13688 17484 13694 17536
rect 14366 17484 14372 17536
rect 14424 17524 14430 17536
rect 14734 17524 14740 17536
rect 14424 17496 14740 17524
rect 14424 17484 14430 17496
rect 14734 17484 14740 17496
rect 14792 17484 14798 17536
rect 16482 17484 16488 17536
rect 16540 17524 16546 17536
rect 17512 17533 17540 17564
rect 17497 17527 17555 17533
rect 17497 17524 17509 17527
rect 16540 17496 17509 17524
rect 16540 17484 16546 17496
rect 17497 17493 17509 17496
rect 17543 17493 17555 17527
rect 17497 17487 17555 17493
rect 18138 17484 18144 17536
rect 18196 17484 18202 17536
rect 18966 17484 18972 17536
rect 19024 17484 19030 17536
rect 19426 17484 19432 17536
rect 19484 17484 19490 17536
rect 1104 17434 23828 17456
rect 1104 17382 2658 17434
rect 2710 17382 2722 17434
rect 2774 17382 2786 17434
rect 2838 17382 2850 17434
rect 2902 17382 2914 17434
rect 2966 17382 2978 17434
rect 3030 17382 8658 17434
rect 8710 17382 8722 17434
rect 8774 17382 8786 17434
rect 8838 17382 8850 17434
rect 8902 17382 8914 17434
rect 8966 17382 8978 17434
rect 9030 17382 14658 17434
rect 14710 17382 14722 17434
rect 14774 17382 14786 17434
rect 14838 17382 14850 17434
rect 14902 17382 14914 17434
rect 14966 17382 14978 17434
rect 15030 17382 20658 17434
rect 20710 17382 20722 17434
rect 20774 17382 20786 17434
rect 20838 17382 20850 17434
rect 20902 17382 20914 17434
rect 20966 17382 20978 17434
rect 21030 17382 23828 17434
rect 1104 17360 23828 17382
rect 4706 17280 4712 17332
rect 4764 17280 4770 17332
rect 6546 17280 6552 17332
rect 6604 17280 6610 17332
rect 6730 17280 6736 17332
rect 6788 17280 6794 17332
rect 6914 17280 6920 17332
rect 6972 17320 6978 17332
rect 9398 17320 9404 17332
rect 6972 17292 8156 17320
rect 6972 17280 6978 17292
rect 4522 17252 4528 17264
rect 3712 17224 4528 17252
rect 1857 17187 1915 17193
rect 1857 17153 1869 17187
rect 1903 17184 1915 17187
rect 3326 17184 3332 17196
rect 1903 17156 3332 17184
rect 1903 17153 1915 17156
rect 1857 17147 1915 17153
rect 3326 17144 3332 17156
rect 3384 17144 3390 17196
rect 3418 17144 3424 17196
rect 3476 17144 3482 17196
rect 3712 17193 3740 17224
rect 4522 17212 4528 17224
rect 4580 17212 4586 17264
rect 6362 17252 6368 17264
rect 4908 17224 6368 17252
rect 3697 17187 3755 17193
rect 3697 17153 3709 17187
rect 3743 17153 3755 17187
rect 3697 17147 3755 17153
rect 3970 17144 3976 17196
rect 4028 17184 4034 17196
rect 4246 17184 4252 17196
rect 4028 17156 4252 17184
rect 4028 17144 4034 17156
rect 4246 17144 4252 17156
rect 4304 17144 4310 17196
rect 4430 17144 4436 17196
rect 4488 17184 4494 17196
rect 4798 17184 4804 17196
rect 4488 17156 4804 17184
rect 4488 17144 4494 17156
rect 4798 17144 4804 17156
rect 4856 17144 4862 17196
rect 934 17076 940 17128
rect 992 17116 998 17128
rect 1581 17119 1639 17125
rect 1581 17116 1593 17119
rect 992 17088 1593 17116
rect 992 17076 998 17088
rect 1581 17085 1593 17088
rect 1627 17085 1639 17119
rect 1581 17079 1639 17085
rect 4157 17119 4215 17125
rect 4157 17085 4169 17119
rect 4203 17116 4215 17119
rect 4908 17116 4936 17224
rect 6362 17212 6368 17224
rect 6420 17212 6426 17264
rect 6564 17252 6592 17280
rect 7469 17255 7527 17261
rect 7469 17252 7481 17255
rect 6564 17224 7481 17252
rect 7469 17221 7481 17224
rect 7515 17221 7527 17255
rect 7469 17215 7527 17221
rect 5074 17193 5080 17196
rect 5068 17147 5080 17193
rect 5074 17144 5080 17147
rect 5132 17144 5138 17196
rect 6457 17187 6515 17193
rect 6457 17184 6469 17187
rect 5828 17156 6469 17184
rect 4203 17088 4936 17116
rect 4203 17085 4215 17088
rect 4157 17079 4215 17085
rect 3605 17051 3663 17057
rect 3605 17017 3617 17051
rect 3651 17048 3663 17051
rect 4614 17048 4620 17060
rect 3651 17020 4620 17048
rect 3651 17017 3663 17020
rect 3605 17011 3663 17017
rect 4614 17008 4620 17020
rect 4672 17008 4678 17060
rect 3050 16940 3056 16992
rect 3108 16980 3114 16992
rect 3237 16983 3295 16989
rect 3237 16980 3249 16983
rect 3108 16952 3249 16980
rect 3108 16940 3114 16952
rect 3237 16949 3249 16952
rect 3283 16949 3295 16983
rect 3237 16943 3295 16949
rect 3881 16983 3939 16989
rect 3881 16949 3893 16983
rect 3927 16980 3939 16983
rect 4246 16980 4252 16992
rect 3927 16952 4252 16980
rect 3927 16949 3939 16952
rect 3881 16943 3939 16949
rect 4246 16940 4252 16952
rect 4304 16940 4310 16992
rect 5166 16940 5172 16992
rect 5224 16980 5230 16992
rect 5828 16980 5856 17156
rect 6457 17153 6469 17156
rect 6503 17153 6515 17187
rect 6457 17147 6515 17153
rect 7098 17116 7104 17128
rect 5920 17088 7104 17116
rect 5920 16992 5948 17088
rect 7098 17076 7104 17088
rect 7156 17076 7162 17128
rect 7285 17119 7343 17125
rect 7285 17085 7297 17119
rect 7331 17116 7343 17119
rect 7484 17116 7512 17215
rect 8128 17184 8156 17292
rect 9140 17292 9404 17320
rect 9140 17184 9168 17292
rect 9398 17280 9404 17292
rect 9456 17320 9462 17332
rect 10873 17323 10931 17329
rect 10873 17320 10885 17323
rect 9456 17292 10885 17320
rect 9456 17280 9462 17292
rect 10873 17289 10885 17292
rect 10919 17289 10931 17323
rect 10873 17283 10931 17289
rect 11517 17323 11575 17329
rect 11517 17289 11529 17323
rect 11563 17289 11575 17323
rect 11517 17283 11575 17289
rect 9217 17255 9275 17261
rect 9217 17221 9229 17255
rect 9263 17252 9275 17255
rect 11532 17252 11560 17283
rect 13262 17280 13268 17332
rect 13320 17280 13326 17332
rect 13630 17280 13636 17332
rect 13688 17280 13694 17332
rect 14737 17323 14795 17329
rect 14737 17289 14749 17323
rect 14783 17320 14795 17323
rect 15654 17320 15660 17332
rect 14783 17292 15660 17320
rect 14783 17289 14795 17292
rect 14737 17283 14795 17289
rect 15654 17280 15660 17292
rect 15712 17280 15718 17332
rect 16393 17323 16451 17329
rect 16393 17289 16405 17323
rect 16439 17320 16451 17323
rect 16850 17320 16856 17332
rect 16439 17292 16856 17320
rect 16439 17289 16451 17292
rect 16393 17283 16451 17289
rect 16850 17280 16856 17292
rect 16908 17280 16914 17332
rect 17034 17280 17040 17332
rect 17092 17320 17098 17332
rect 17862 17320 17868 17332
rect 17092 17292 17868 17320
rect 17092 17280 17098 17292
rect 17862 17280 17868 17292
rect 17920 17320 17926 17332
rect 17957 17323 18015 17329
rect 17957 17320 17969 17323
rect 17920 17292 17969 17320
rect 17920 17280 17926 17292
rect 17957 17289 17969 17292
rect 18003 17289 18015 17323
rect 17957 17283 18015 17289
rect 18138 17280 18144 17332
rect 18196 17280 18202 17332
rect 18966 17280 18972 17332
rect 19024 17280 19030 17332
rect 9263 17224 11560 17252
rect 12152 17255 12210 17261
rect 9263 17221 9275 17224
rect 9217 17215 9275 17221
rect 12152 17221 12164 17255
rect 12198 17252 12210 17255
rect 13170 17252 13176 17264
rect 12198 17224 13176 17252
rect 12198 17221 12210 17224
rect 12152 17215 12210 17221
rect 13170 17212 13176 17224
rect 13228 17212 13234 17264
rect 13648 17252 13676 17280
rect 13372 17224 13676 17252
rect 9309 17187 9367 17193
rect 9309 17184 9321 17187
rect 8128 17156 9321 17184
rect 9309 17153 9321 17156
rect 9355 17153 9367 17187
rect 9309 17147 9367 17153
rect 9585 17187 9643 17193
rect 9585 17153 9597 17187
rect 9631 17153 9643 17187
rect 9585 17147 9643 17153
rect 9600 17116 9628 17147
rect 11422 17144 11428 17196
rect 11480 17144 11486 17196
rect 11698 17144 11704 17196
rect 11756 17144 11762 17196
rect 13372 17193 13400 17224
rect 14366 17212 14372 17264
rect 14424 17212 14430 17264
rect 18156 17252 18184 17280
rect 15028 17224 18184 17252
rect 18984 17252 19012 17280
rect 18984 17224 20024 17252
rect 13357 17187 13415 17193
rect 13357 17153 13369 17187
rect 13403 17153 13415 17187
rect 13357 17147 13415 17153
rect 13624 17187 13682 17193
rect 13624 17153 13636 17187
rect 13670 17184 13682 17187
rect 14384 17184 14412 17212
rect 15028 17193 15056 17224
rect 15286 17193 15292 17196
rect 13670 17156 14412 17184
rect 15013 17187 15071 17193
rect 13670 17153 13682 17156
rect 13624 17147 13682 17153
rect 15013 17153 15025 17187
rect 15059 17153 15071 17187
rect 15280 17184 15292 17193
rect 15247 17156 15292 17184
rect 15013 17147 15071 17153
rect 15280 17147 15292 17156
rect 15286 17144 15292 17147
rect 15344 17144 15350 17196
rect 16669 17187 16727 17193
rect 16669 17153 16681 17187
rect 16715 17184 16727 17187
rect 16850 17184 16856 17196
rect 16715 17156 16856 17184
rect 16715 17153 16727 17156
rect 16669 17147 16727 17153
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 19610 17144 19616 17196
rect 19668 17193 19674 17196
rect 19996 17193 20024 17224
rect 19668 17147 19680 17193
rect 19981 17187 20039 17193
rect 19981 17153 19993 17187
rect 20027 17153 20039 17187
rect 19981 17147 20039 17153
rect 20248 17187 20306 17193
rect 20248 17153 20260 17187
rect 20294 17184 20306 17187
rect 21174 17184 21180 17196
rect 20294 17156 21180 17184
rect 20294 17153 20306 17156
rect 20248 17147 20306 17153
rect 19668 17144 19674 17147
rect 21174 17144 21180 17156
rect 21232 17144 21238 17196
rect 23017 17187 23075 17193
rect 23017 17184 23029 17187
rect 22066 17156 23029 17184
rect 7331 17088 7420 17116
rect 7484 17088 9628 17116
rect 11440 17116 11468 17144
rect 11885 17119 11943 17125
rect 11885 17116 11897 17119
rect 11440 17088 11897 17116
rect 7331 17085 7343 17088
rect 7285 17079 7343 17085
rect 6549 17051 6607 17057
rect 6549 17017 6561 17051
rect 6595 17048 6607 17051
rect 7006 17048 7012 17060
rect 6595 17020 7012 17048
rect 6595 17017 6607 17020
rect 6549 17011 6607 17017
rect 7006 17008 7012 17020
rect 7064 17008 7070 17060
rect 7392 17048 7420 17088
rect 11885 17085 11897 17088
rect 11931 17085 11943 17119
rect 11885 17079 11943 17085
rect 19889 17119 19947 17125
rect 19889 17085 19901 17119
rect 19935 17085 19947 17119
rect 19889 17079 19947 17085
rect 11514 17048 11520 17060
rect 7392 17020 11520 17048
rect 11514 17008 11520 17020
rect 11572 17008 11578 17060
rect 5224 16952 5856 16980
rect 5224 16940 5230 16952
rect 5902 16940 5908 16992
rect 5960 16940 5966 16992
rect 6181 16983 6239 16989
rect 6181 16949 6193 16983
rect 6227 16980 6239 16983
rect 6454 16980 6460 16992
rect 6227 16952 6460 16980
rect 6227 16949 6239 16952
rect 6181 16943 6239 16949
rect 6454 16940 6460 16952
rect 6512 16940 6518 16992
rect 9401 16983 9459 16989
rect 9401 16949 9413 16983
rect 9447 16980 9459 16983
rect 10502 16980 10508 16992
rect 9447 16952 10508 16980
rect 9447 16949 9459 16952
rect 9401 16943 9459 16949
rect 10502 16940 10508 16952
rect 10560 16940 10566 16992
rect 18506 16940 18512 16992
rect 18564 16940 18570 16992
rect 19518 16940 19524 16992
rect 19576 16980 19582 16992
rect 19904 16980 19932 17079
rect 21361 17051 21419 17057
rect 21361 17017 21373 17051
rect 21407 17048 21419 17051
rect 22066 17048 22094 17156
rect 23017 17153 23029 17156
rect 23063 17153 23075 17187
rect 23017 17147 23075 17153
rect 23290 17076 23296 17128
rect 23348 17076 23354 17128
rect 21407 17020 22094 17048
rect 21407 17017 21419 17020
rect 21361 17011 21419 17017
rect 21082 16980 21088 16992
rect 19576 16952 21088 16980
rect 19576 16940 19582 16952
rect 21082 16940 21088 16952
rect 21140 16940 21146 16992
rect 1104 16890 23828 16912
rect 1104 16838 1918 16890
rect 1970 16838 1982 16890
rect 2034 16838 2046 16890
rect 2098 16838 2110 16890
rect 2162 16838 2174 16890
rect 2226 16838 2238 16890
rect 2290 16838 7918 16890
rect 7970 16838 7982 16890
rect 8034 16838 8046 16890
rect 8098 16838 8110 16890
rect 8162 16838 8174 16890
rect 8226 16838 8238 16890
rect 8290 16838 13918 16890
rect 13970 16838 13982 16890
rect 14034 16838 14046 16890
rect 14098 16838 14110 16890
rect 14162 16838 14174 16890
rect 14226 16838 14238 16890
rect 14290 16838 19918 16890
rect 19970 16838 19982 16890
rect 20034 16838 20046 16890
rect 20098 16838 20110 16890
rect 20162 16838 20174 16890
rect 20226 16838 20238 16890
rect 20290 16838 23828 16890
rect 1104 16816 23828 16838
rect 6086 16776 6092 16788
rect 3068 16748 6092 16776
rect 3068 16649 3096 16748
rect 6086 16736 6092 16748
rect 6144 16736 6150 16788
rect 6178 16736 6184 16788
rect 6236 16776 6242 16788
rect 6733 16779 6791 16785
rect 6733 16776 6745 16779
rect 6236 16748 6745 16776
rect 6236 16736 6242 16748
rect 6733 16745 6745 16748
rect 6779 16745 6791 16779
rect 6733 16739 6791 16745
rect 6822 16736 6828 16788
rect 6880 16736 6886 16788
rect 11606 16736 11612 16788
rect 11664 16736 11670 16788
rect 18414 16736 18420 16788
rect 18472 16776 18478 16788
rect 19886 16776 19892 16788
rect 18472 16748 19892 16776
rect 18472 16736 18478 16748
rect 19886 16736 19892 16748
rect 19944 16736 19950 16788
rect 21174 16736 21180 16788
rect 21232 16736 21238 16788
rect 3053 16643 3111 16649
rect 3053 16609 3065 16643
rect 3099 16609 3111 16643
rect 3053 16603 3111 16609
rect 3234 16600 3240 16652
rect 3292 16640 3298 16652
rect 5166 16640 5172 16652
rect 3292 16612 5172 16640
rect 3292 16600 3298 16612
rect 2130 16532 2136 16584
rect 2188 16532 2194 16584
rect 3988 16581 4016 16612
rect 5166 16600 5172 16612
rect 5224 16600 5230 16652
rect 6365 16643 6423 16649
rect 6365 16609 6377 16643
rect 6411 16640 6423 16643
rect 6840 16640 6868 16736
rect 8389 16711 8447 16717
rect 8389 16677 8401 16711
rect 8435 16677 8447 16711
rect 8389 16671 8447 16677
rect 8404 16640 8432 16671
rect 9030 16668 9036 16720
rect 9088 16668 9094 16720
rect 12345 16711 12403 16717
rect 12345 16708 12357 16711
rect 12268 16680 12357 16708
rect 12268 16649 12296 16680
rect 12345 16677 12357 16680
rect 12391 16677 12403 16711
rect 18693 16711 18751 16717
rect 12345 16671 12403 16677
rect 18064 16680 18644 16708
rect 18064 16652 18092 16680
rect 6411 16612 6868 16640
rect 6932 16612 8432 16640
rect 12253 16643 12311 16649
rect 6411 16609 6423 16612
rect 6365 16603 6423 16609
rect 2685 16575 2743 16581
rect 2685 16572 2697 16575
rect 2424 16544 2697 16572
rect 2424 16448 2452 16544
rect 2685 16541 2697 16544
rect 2731 16541 2743 16575
rect 2685 16535 2743 16541
rect 3973 16575 4031 16581
rect 3973 16541 3985 16575
rect 4019 16541 4031 16575
rect 3973 16535 4031 16541
rect 4341 16575 4399 16581
rect 4341 16541 4353 16575
rect 4387 16572 4399 16575
rect 5810 16572 5816 16584
rect 4387 16544 5816 16572
rect 4387 16541 4399 16544
rect 4341 16535 4399 16541
rect 5810 16532 5816 16544
rect 5868 16532 5874 16584
rect 6109 16575 6167 16581
rect 6109 16541 6121 16575
rect 6155 16572 6167 16575
rect 6270 16572 6276 16584
rect 6155 16544 6276 16572
rect 6155 16541 6167 16544
rect 6109 16535 6167 16541
rect 6270 16532 6276 16544
rect 6328 16532 6334 16584
rect 6932 16572 6960 16612
rect 12253 16609 12265 16643
rect 12299 16609 12311 16643
rect 12253 16603 12311 16609
rect 13725 16643 13783 16649
rect 13725 16609 13737 16643
rect 13771 16640 13783 16643
rect 14366 16640 14372 16652
rect 13771 16612 14372 16640
rect 13771 16609 13783 16612
rect 13725 16603 13783 16609
rect 14366 16600 14372 16612
rect 14424 16600 14430 16652
rect 17681 16643 17739 16649
rect 17681 16609 17693 16643
rect 17727 16640 17739 16643
rect 18046 16640 18052 16652
rect 17727 16612 18052 16640
rect 17727 16609 17739 16612
rect 17681 16603 17739 16609
rect 18046 16600 18052 16612
rect 18104 16600 18110 16652
rect 18616 16640 18644 16680
rect 18693 16677 18705 16711
rect 18739 16708 18751 16711
rect 19794 16708 19800 16720
rect 18739 16680 19800 16708
rect 18739 16677 18751 16680
rect 18693 16671 18751 16677
rect 19794 16668 19800 16680
rect 19852 16668 19858 16720
rect 21726 16668 21732 16720
rect 21784 16668 21790 16720
rect 18616 16612 19288 16640
rect 11333 16575 11391 16581
rect 11333 16572 11345 16575
rect 6656 16544 6960 16572
rect 8220 16544 11345 16572
rect 2777 16507 2835 16513
rect 2777 16473 2789 16507
rect 2823 16504 2835 16507
rect 4154 16504 4160 16516
rect 2823 16476 4160 16504
rect 2823 16473 2835 16476
rect 2777 16467 2835 16473
rect 4154 16464 4160 16476
rect 4212 16464 4218 16516
rect 4893 16507 4951 16513
rect 4893 16473 4905 16507
rect 4939 16504 4951 16507
rect 6656 16504 6684 16544
rect 8220 16513 8248 16544
rect 11333 16541 11345 16544
rect 11379 16541 11391 16575
rect 11333 16535 11391 16541
rect 13458 16575 13516 16581
rect 13458 16541 13470 16575
rect 13504 16541 13516 16575
rect 15838 16572 15844 16584
rect 13458 16535 13516 16541
rect 13639 16544 15844 16572
rect 8205 16507 8263 16513
rect 8205 16504 8217 16507
rect 4939 16476 5856 16504
rect 4939 16473 4951 16476
rect 4893 16467 4951 16473
rect 1210 16396 1216 16448
rect 1268 16436 1274 16448
rect 2041 16439 2099 16445
rect 2041 16436 2053 16439
rect 1268 16408 2053 16436
rect 1268 16396 1274 16408
rect 2041 16405 2053 16408
rect 2087 16405 2099 16439
rect 2041 16399 2099 16405
rect 2406 16396 2412 16448
rect 2464 16396 2470 16448
rect 3418 16396 3424 16448
rect 3476 16436 3482 16448
rect 3605 16439 3663 16445
rect 3605 16436 3617 16439
rect 3476 16408 3617 16436
rect 3476 16396 3482 16408
rect 3605 16405 3617 16408
rect 3651 16405 3663 16439
rect 3605 16399 3663 16405
rect 4062 16396 4068 16448
rect 4120 16396 4126 16448
rect 4985 16439 5043 16445
rect 4985 16405 4997 16439
rect 5031 16436 5043 16439
rect 5442 16436 5448 16448
rect 5031 16408 5448 16436
rect 5031 16405 5043 16408
rect 4985 16399 5043 16405
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 5828 16436 5856 16476
rect 6104 16476 6684 16504
rect 7760 16476 8217 16504
rect 6104 16436 6132 16476
rect 7760 16448 7788 16476
rect 8205 16473 8217 16476
rect 8251 16473 8263 16507
rect 8205 16467 8263 16473
rect 8662 16464 8668 16516
rect 8720 16464 8726 16516
rect 8757 16507 8815 16513
rect 8757 16473 8769 16507
rect 8803 16504 8815 16507
rect 9398 16504 9404 16516
rect 8803 16476 9404 16504
rect 8803 16473 8815 16476
rect 8757 16467 8815 16473
rect 9398 16464 9404 16476
rect 9456 16464 9462 16516
rect 5828 16408 6132 16436
rect 7742 16396 7748 16448
rect 7800 16396 7806 16448
rect 8294 16396 8300 16448
rect 8352 16396 8358 16448
rect 8680 16436 8708 16464
rect 8941 16439 8999 16445
rect 8941 16436 8953 16439
rect 8680 16408 8953 16436
rect 8941 16405 8953 16408
rect 8987 16405 8999 16439
rect 8941 16399 8999 16405
rect 9858 16396 9864 16448
rect 9916 16396 9922 16448
rect 11348 16436 11376 16535
rect 13464 16504 13492 16535
rect 13538 16504 13544 16516
rect 13464 16476 13544 16504
rect 13538 16464 13544 16476
rect 13596 16464 13602 16516
rect 13170 16436 13176 16448
rect 11348 16408 13176 16436
rect 13170 16396 13176 16408
rect 13228 16436 13234 16448
rect 13639 16436 13667 16544
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 18414 16532 18420 16584
rect 18472 16532 18478 16584
rect 19260 16581 19288 16612
rect 21082 16600 21088 16652
rect 21140 16640 21146 16652
rect 21744 16640 21772 16668
rect 21140 16612 21772 16640
rect 21140 16600 21146 16612
rect 22186 16600 22192 16652
rect 22244 16640 22250 16652
rect 22465 16643 22523 16649
rect 22465 16640 22477 16643
rect 22244 16612 22477 16640
rect 22244 16600 22250 16612
rect 22465 16609 22477 16612
rect 22511 16609 22523 16643
rect 22465 16603 22523 16609
rect 19245 16575 19303 16581
rect 19245 16541 19257 16575
rect 19291 16541 19303 16575
rect 19245 16535 19303 16541
rect 21729 16575 21787 16581
rect 21729 16541 21741 16575
rect 21775 16541 21787 16575
rect 21729 16535 21787 16541
rect 22833 16575 22891 16581
rect 22833 16541 22845 16575
rect 22879 16541 22891 16575
rect 22833 16535 22891 16541
rect 14093 16507 14151 16513
rect 14093 16504 14105 16507
rect 13832 16476 14105 16504
rect 13832 16448 13860 16476
rect 14093 16473 14105 16476
rect 14139 16473 14151 16507
rect 14093 16467 14151 16473
rect 15930 16464 15936 16516
rect 15988 16464 15994 16516
rect 18598 16464 18604 16516
rect 18656 16504 18662 16516
rect 18969 16507 19027 16513
rect 18969 16504 18981 16507
rect 18656 16476 18981 16504
rect 18656 16464 18662 16476
rect 18969 16473 18981 16476
rect 19015 16473 19027 16507
rect 20818 16507 20876 16513
rect 20818 16504 20830 16507
rect 18969 16467 19027 16473
rect 19260 16476 20830 16504
rect 19260 16448 19288 16476
rect 20818 16473 20830 16476
rect 20864 16504 20876 16507
rect 21744 16504 21772 16535
rect 20864 16476 21772 16504
rect 22848 16504 22876 16535
rect 23014 16532 23020 16584
rect 23072 16532 23078 16584
rect 22848 16476 23152 16504
rect 20864 16473 20876 16476
rect 20818 16467 20876 16473
rect 23124 16448 23152 16476
rect 23198 16464 23204 16516
rect 23256 16504 23262 16516
rect 23293 16507 23351 16513
rect 23293 16504 23305 16507
rect 23256 16476 23305 16504
rect 23256 16464 23262 16476
rect 23293 16473 23305 16476
rect 23339 16473 23351 16507
rect 23293 16467 23351 16473
rect 13228 16408 13667 16436
rect 13228 16396 13234 16408
rect 13814 16396 13820 16448
rect 13872 16396 13878 16448
rect 16206 16396 16212 16448
rect 16264 16436 16270 16448
rect 17773 16439 17831 16445
rect 17773 16436 17785 16439
rect 16264 16408 17785 16436
rect 16264 16396 16270 16408
rect 17773 16405 17785 16408
rect 17819 16405 17831 16439
rect 17773 16399 17831 16405
rect 18230 16396 18236 16448
rect 18288 16436 18294 16448
rect 18509 16439 18567 16445
rect 18509 16436 18521 16439
rect 18288 16408 18521 16436
rect 18288 16396 18294 16408
rect 18509 16405 18521 16408
rect 18555 16405 18567 16439
rect 18509 16399 18567 16405
rect 19242 16396 19248 16448
rect 19300 16396 19306 16448
rect 19334 16396 19340 16448
rect 19392 16396 19398 16448
rect 19702 16396 19708 16448
rect 19760 16396 19766 16448
rect 21910 16396 21916 16448
rect 21968 16396 21974 16448
rect 22738 16396 22744 16448
rect 22796 16396 22802 16448
rect 23106 16396 23112 16448
rect 23164 16396 23170 16448
rect 1104 16346 23828 16368
rect 1104 16294 2658 16346
rect 2710 16294 2722 16346
rect 2774 16294 2786 16346
rect 2838 16294 2850 16346
rect 2902 16294 2914 16346
rect 2966 16294 2978 16346
rect 3030 16294 8658 16346
rect 8710 16294 8722 16346
rect 8774 16294 8786 16346
rect 8838 16294 8850 16346
rect 8902 16294 8914 16346
rect 8966 16294 8978 16346
rect 9030 16294 14658 16346
rect 14710 16294 14722 16346
rect 14774 16294 14786 16346
rect 14838 16294 14850 16346
rect 14902 16294 14914 16346
rect 14966 16294 14978 16346
rect 15030 16294 20658 16346
rect 20710 16294 20722 16346
rect 20774 16294 20786 16346
rect 20838 16294 20850 16346
rect 20902 16294 20914 16346
rect 20966 16294 20978 16346
rect 21030 16294 23828 16346
rect 1104 16272 23828 16294
rect 3326 16192 3332 16244
rect 3384 16192 3390 16244
rect 3694 16192 3700 16244
rect 3752 16232 3758 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 3752 16204 6193 16232
rect 3752 16192 3758 16204
rect 6181 16201 6193 16204
rect 6227 16201 6239 16235
rect 6181 16195 6239 16201
rect 6549 16235 6607 16241
rect 6549 16201 6561 16235
rect 6595 16232 6607 16235
rect 9766 16232 9772 16244
rect 6595 16204 9772 16232
rect 6595 16201 6607 16204
rect 6549 16195 6607 16201
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 11514 16192 11520 16244
rect 11572 16192 11578 16244
rect 12066 16192 12072 16244
rect 12124 16192 12130 16244
rect 13262 16232 13268 16244
rect 13188 16204 13268 16232
rect 1486 16124 1492 16176
rect 1544 16164 1550 16176
rect 1544 16136 2360 16164
rect 1544 16124 1550 16136
rect 1854 16056 1860 16108
rect 1912 16056 1918 16108
rect 2332 16105 2360 16136
rect 3418 16124 3424 16176
rect 3476 16164 3482 16176
rect 3476 16136 4016 16164
rect 3476 16124 3482 16136
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16065 2099 16099
rect 2041 16059 2099 16065
rect 2317 16099 2375 16105
rect 2317 16065 2329 16099
rect 2363 16096 2375 16099
rect 2685 16099 2743 16105
rect 2363 16068 2636 16096
rect 2363 16065 2375 16068
rect 2317 16059 2375 16065
rect 934 15988 940 16040
rect 992 16028 998 16040
rect 1581 16031 1639 16037
rect 1581 16028 1593 16031
rect 992 16000 1593 16028
rect 992 15988 998 16000
rect 1581 15997 1593 16000
rect 1627 15997 1639 16031
rect 1581 15991 1639 15997
rect 1670 15988 1676 16040
rect 1728 16028 1734 16040
rect 2056 16028 2084 16059
rect 1728 16000 2084 16028
rect 2133 16031 2191 16037
rect 1728 15988 1734 16000
rect 2133 15997 2145 16031
rect 2179 16028 2191 16031
rect 2498 16028 2504 16040
rect 2179 16000 2504 16028
rect 2179 15997 2191 16000
rect 2133 15991 2191 15997
rect 2498 15988 2504 16000
rect 2556 15988 2562 16040
rect 2608 16028 2636 16068
rect 2685 16065 2697 16099
rect 2731 16096 2743 16099
rect 3694 16096 3700 16108
rect 2731 16068 3700 16096
rect 2731 16065 2743 16068
rect 2685 16059 2743 16065
rect 3694 16056 3700 16068
rect 3752 16056 3758 16108
rect 3988 16096 4016 16136
rect 4062 16124 4068 16176
rect 4120 16164 4126 16176
rect 4120 16136 4844 16164
rect 4120 16124 4126 16136
rect 4816 16105 4844 16136
rect 4890 16124 4896 16176
rect 4948 16164 4954 16176
rect 5046 16167 5104 16173
rect 5046 16164 5058 16167
rect 4948 16136 5058 16164
rect 4948 16124 4954 16136
rect 5046 16133 5058 16136
rect 5092 16133 5104 16167
rect 10597 16167 10655 16173
rect 5046 16127 5104 16133
rect 7024 16136 8156 16164
rect 7024 16108 7052 16136
rect 4442 16099 4500 16105
rect 4442 16096 4454 16099
rect 3988 16068 4454 16096
rect 4442 16065 4454 16068
rect 4488 16065 4500 16099
rect 4442 16059 4500 16065
rect 4801 16099 4859 16105
rect 4801 16065 4813 16099
rect 4847 16065 4859 16099
rect 4801 16059 4859 16065
rect 6638 16056 6644 16108
rect 6696 16056 6702 16108
rect 7006 16056 7012 16108
rect 7064 16056 7070 16108
rect 7834 16056 7840 16108
rect 7892 16105 7898 16108
rect 8128 16105 8156 16136
rect 10597 16133 10609 16167
rect 10643 16164 10655 16167
rect 11882 16164 11888 16176
rect 10643 16136 11888 16164
rect 10643 16133 10655 16136
rect 10597 16127 10655 16133
rect 11882 16124 11888 16136
rect 11940 16164 11946 16176
rect 13188 16173 13216 16204
rect 13262 16192 13268 16204
rect 13320 16192 13326 16244
rect 14366 16192 14372 16244
rect 14424 16192 14430 16244
rect 15838 16192 15844 16244
rect 15896 16232 15902 16244
rect 15896 16204 16988 16232
rect 15896 16192 15902 16204
rect 11977 16167 12035 16173
rect 11977 16164 11989 16167
rect 11940 16136 11989 16164
rect 11940 16124 11946 16136
rect 11977 16133 11989 16136
rect 12023 16133 12035 16167
rect 11977 16127 12035 16133
rect 13182 16167 13240 16173
rect 13182 16133 13194 16167
rect 13228 16133 13240 16167
rect 13182 16127 13240 16133
rect 13906 16124 13912 16176
rect 13964 16164 13970 16176
rect 16960 16173 16988 16204
rect 17034 16192 17040 16244
rect 17092 16232 17098 16244
rect 18417 16235 18475 16241
rect 18417 16232 18429 16235
rect 17092 16204 18429 16232
rect 17092 16192 17098 16204
rect 18417 16201 18429 16204
rect 18463 16232 18475 16235
rect 19518 16232 19524 16244
rect 18463 16204 19524 16232
rect 18463 16201 18475 16204
rect 18417 16195 18475 16201
rect 19518 16192 19524 16204
rect 19576 16192 19582 16244
rect 19794 16192 19800 16244
rect 19852 16232 19858 16244
rect 20625 16235 20683 16241
rect 20625 16232 20637 16235
rect 19852 16204 20637 16232
rect 19852 16192 19858 16204
rect 20625 16201 20637 16204
rect 20671 16201 20683 16235
rect 20625 16195 20683 16201
rect 16945 16167 17003 16173
rect 13964 16136 16252 16164
rect 13964 16124 13970 16136
rect 7892 16096 7904 16105
rect 8113 16099 8171 16105
rect 7892 16068 7937 16096
rect 7892 16059 7904 16068
rect 8113 16065 8125 16099
rect 8159 16065 8171 16099
rect 8113 16059 8171 16065
rect 8205 16099 8263 16105
rect 8205 16065 8217 16099
rect 8251 16065 8263 16099
rect 8205 16059 8263 16065
rect 13449 16099 13507 16105
rect 13449 16065 13461 16099
rect 13495 16096 13507 16099
rect 13814 16096 13820 16108
rect 13495 16068 13820 16096
rect 13495 16065 13507 16068
rect 13449 16059 13507 16065
rect 7892 16056 7898 16059
rect 3602 16028 3608 16040
rect 2608 16000 3608 16028
rect 3602 15988 3608 16000
rect 3660 15988 3666 16040
rect 4706 15988 4712 16040
rect 4764 15988 4770 16040
rect 7006 15960 7012 15972
rect 6104 15932 7012 15960
rect 2498 15852 2504 15904
rect 2556 15852 2562 15904
rect 3237 15895 3295 15901
rect 3237 15861 3249 15895
rect 3283 15892 3295 15895
rect 3694 15892 3700 15904
rect 3283 15864 3700 15892
rect 3283 15861 3295 15864
rect 3237 15855 3295 15861
rect 3694 15852 3700 15864
rect 3752 15852 3758 15904
rect 4522 15852 4528 15904
rect 4580 15892 4586 15904
rect 6104 15892 6132 15932
rect 7006 15920 7012 15932
rect 7064 15920 7070 15972
rect 4580 15864 6132 15892
rect 4580 15852 4586 15864
rect 6362 15852 6368 15904
rect 6420 15892 6426 15904
rect 6733 15895 6791 15901
rect 6733 15892 6745 15895
rect 6420 15864 6745 15892
rect 6420 15852 6426 15864
rect 6733 15861 6745 15864
rect 6779 15861 6791 15895
rect 6733 15855 6791 15861
rect 6822 15852 6828 15904
rect 6880 15892 6886 15904
rect 8220 15892 8248 16059
rect 13814 16056 13820 16068
rect 13872 16096 13878 16108
rect 13872 16068 14228 16096
rect 13872 16056 13878 16068
rect 11330 15988 11336 16040
rect 11388 15988 11394 16040
rect 13722 15988 13728 16040
rect 13780 16028 13786 16040
rect 14093 16031 14151 16037
rect 14093 16028 14105 16031
rect 13780 16000 14105 16028
rect 13780 15988 13786 16000
rect 14093 15997 14105 16000
rect 14139 15997 14151 16031
rect 14200 16028 14228 16068
rect 14366 16056 14372 16108
rect 14424 16096 14430 16108
rect 14461 16099 14519 16105
rect 14461 16096 14473 16099
rect 14424 16068 14473 16096
rect 14424 16056 14430 16068
rect 14461 16065 14473 16068
rect 14507 16096 14519 16099
rect 14550 16096 14556 16108
rect 14507 16068 14556 16096
rect 14507 16065 14519 16068
rect 14461 16059 14519 16065
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 15004 16099 15062 16105
rect 15004 16065 15016 16099
rect 15050 16096 15062 16099
rect 15286 16096 15292 16108
rect 15050 16068 15292 16096
rect 15050 16065 15062 16068
rect 15004 16059 15062 16065
rect 15286 16056 15292 16068
rect 15344 16056 15350 16108
rect 16224 16105 16252 16136
rect 16945 16133 16957 16167
rect 16991 16133 17003 16167
rect 16945 16127 17003 16133
rect 17862 16124 17868 16176
rect 17920 16164 17926 16176
rect 18785 16167 18843 16173
rect 18785 16164 18797 16167
rect 17920 16136 18797 16164
rect 17920 16124 17926 16136
rect 18785 16133 18797 16136
rect 18831 16133 18843 16167
rect 23106 16164 23112 16176
rect 18785 16127 18843 16133
rect 21560 16136 23112 16164
rect 16209 16099 16267 16105
rect 16209 16065 16221 16099
rect 16255 16065 16267 16099
rect 16209 16059 16267 16065
rect 14737 16031 14795 16037
rect 14737 16028 14749 16031
rect 14200 16000 14749 16028
rect 14093 15991 14151 15997
rect 14737 15997 14749 16000
rect 14783 15997 14795 16031
rect 14737 15991 14795 15997
rect 9490 15920 9496 15972
rect 9548 15920 9554 15972
rect 10321 15963 10379 15969
rect 10321 15929 10333 15963
rect 10367 15960 10379 15963
rect 10689 15963 10747 15969
rect 10689 15960 10701 15963
rect 10367 15932 10701 15960
rect 10367 15929 10379 15932
rect 10321 15923 10379 15929
rect 10689 15929 10701 15932
rect 10735 15929 10747 15963
rect 10689 15923 10747 15929
rect 11701 15963 11759 15969
rect 11701 15929 11713 15963
rect 11747 15960 11759 15963
rect 11790 15960 11796 15972
rect 11747 15932 11796 15960
rect 11747 15929 11759 15932
rect 11701 15923 11759 15929
rect 11790 15920 11796 15932
rect 11848 15920 11854 15972
rect 6880 15864 8248 15892
rect 6880 15852 6886 15864
rect 9674 15852 9680 15904
rect 9732 15892 9738 15904
rect 10137 15895 10195 15901
rect 10137 15892 10149 15895
rect 9732 15864 10149 15892
rect 9732 15852 9738 15864
rect 10137 15861 10149 15864
rect 10183 15861 10195 15895
rect 10137 15855 10195 15861
rect 13446 15852 13452 15904
rect 13504 15892 13510 15904
rect 13541 15895 13599 15901
rect 13541 15892 13553 15895
rect 13504 15864 13553 15892
rect 13504 15852 13510 15864
rect 13541 15861 13553 15864
rect 13587 15861 13599 15895
rect 14752 15892 14780 15991
rect 16224 15960 16252 16059
rect 16666 16056 16672 16108
rect 16724 16056 16730 16108
rect 21560 16105 21588 16136
rect 23106 16124 23112 16136
rect 23164 16124 23170 16176
rect 21545 16099 21603 16105
rect 21545 16065 21557 16099
rect 21591 16065 21603 16099
rect 21545 16059 21603 16065
rect 22002 16056 22008 16108
rect 22060 16056 22066 16108
rect 20346 15988 20352 16040
rect 20404 16028 20410 16040
rect 21177 16031 21235 16037
rect 21177 16028 21189 16031
rect 20404 16000 21189 16028
rect 20404 15988 20410 16000
rect 21177 15997 21189 16000
rect 21223 15997 21235 16031
rect 21177 15991 21235 15997
rect 22094 15988 22100 16040
rect 22152 15988 22158 16040
rect 22922 15988 22928 16040
rect 22980 16028 22986 16040
rect 23385 16031 23443 16037
rect 23385 16028 23397 16031
rect 22980 16000 23397 16028
rect 22980 15988 22986 16000
rect 23385 15997 23397 16000
rect 23431 15997 23443 16031
rect 23385 15991 23443 15997
rect 19058 15960 19064 15972
rect 16224 15932 19064 15960
rect 19058 15920 19064 15932
rect 19116 15960 19122 15972
rect 20073 15963 20131 15969
rect 20073 15960 20085 15963
rect 19116 15932 20085 15960
rect 19116 15920 19122 15932
rect 20073 15929 20085 15932
rect 20119 15960 20131 15963
rect 21634 15960 21640 15972
rect 20119 15932 21640 15960
rect 20119 15929 20131 15932
rect 20073 15923 20131 15929
rect 21634 15920 21640 15932
rect 21692 15920 21698 15972
rect 21913 15963 21971 15969
rect 21913 15929 21925 15963
rect 21959 15960 21971 15963
rect 23198 15960 23204 15972
rect 21959 15932 23204 15960
rect 21959 15929 21971 15932
rect 21913 15923 21971 15929
rect 23198 15920 23204 15932
rect 23256 15920 23262 15972
rect 15102 15892 15108 15904
rect 14752 15864 15108 15892
rect 13541 15855 13599 15861
rect 15102 15852 15108 15864
rect 15160 15852 15166 15904
rect 16114 15852 16120 15904
rect 16172 15852 16178 15904
rect 16301 15895 16359 15901
rect 16301 15861 16313 15895
rect 16347 15892 16359 15895
rect 16574 15892 16580 15904
rect 16347 15864 16580 15892
rect 16347 15861 16359 15864
rect 16301 15855 16359 15861
rect 16574 15852 16580 15864
rect 16632 15852 16638 15904
rect 16761 15895 16819 15901
rect 16761 15861 16773 15895
rect 16807 15892 16819 15895
rect 17954 15892 17960 15904
rect 16807 15864 17960 15892
rect 16807 15861 16819 15864
rect 16761 15855 16819 15861
rect 17954 15852 17960 15864
rect 18012 15852 18018 15904
rect 21450 15852 21456 15904
rect 21508 15852 21514 15904
rect 22554 15852 22560 15904
rect 22612 15892 22618 15904
rect 22741 15895 22799 15901
rect 22741 15892 22753 15895
rect 22612 15864 22753 15892
rect 22612 15852 22618 15864
rect 22741 15861 22753 15864
rect 22787 15861 22799 15895
rect 22741 15855 22799 15861
rect 22830 15852 22836 15904
rect 22888 15852 22894 15904
rect 1104 15802 23828 15824
rect 1104 15750 1918 15802
rect 1970 15750 1982 15802
rect 2034 15750 2046 15802
rect 2098 15750 2110 15802
rect 2162 15750 2174 15802
rect 2226 15750 2238 15802
rect 2290 15750 7918 15802
rect 7970 15750 7982 15802
rect 8034 15750 8046 15802
rect 8098 15750 8110 15802
rect 8162 15750 8174 15802
rect 8226 15750 8238 15802
rect 8290 15750 13918 15802
rect 13970 15750 13982 15802
rect 14034 15750 14046 15802
rect 14098 15750 14110 15802
rect 14162 15750 14174 15802
rect 14226 15750 14238 15802
rect 14290 15750 19918 15802
rect 19970 15750 19982 15802
rect 20034 15750 20046 15802
rect 20098 15750 20110 15802
rect 20162 15750 20174 15802
rect 20226 15750 20238 15802
rect 20290 15750 23828 15802
rect 1104 15728 23828 15750
rect 1673 15691 1731 15697
rect 1673 15657 1685 15691
rect 1719 15688 1731 15691
rect 3605 15691 3663 15697
rect 1719 15660 3464 15688
rect 1719 15657 1731 15660
rect 1673 15651 1731 15657
rect 3436 15620 3464 15660
rect 3605 15657 3617 15691
rect 3651 15688 3663 15691
rect 3878 15688 3884 15700
rect 3651 15660 3884 15688
rect 3651 15657 3663 15660
rect 3605 15651 3663 15657
rect 3878 15648 3884 15660
rect 3936 15648 3942 15700
rect 3973 15691 4031 15697
rect 3973 15657 3985 15691
rect 4019 15688 4031 15691
rect 4706 15688 4712 15700
rect 4019 15660 4712 15688
rect 4019 15657 4031 15660
rect 3973 15651 4031 15657
rect 4706 15648 4712 15660
rect 4764 15648 4770 15700
rect 4798 15648 4804 15700
rect 4856 15688 4862 15700
rect 7285 15691 7343 15697
rect 7285 15688 7297 15691
rect 4856 15660 7297 15688
rect 4856 15648 4862 15660
rect 7285 15657 7297 15660
rect 7331 15657 7343 15691
rect 7285 15651 7343 15657
rect 7377 15691 7435 15697
rect 7377 15657 7389 15691
rect 7423 15688 7435 15691
rect 7466 15688 7472 15700
rect 7423 15660 7472 15688
rect 7423 15657 7435 15660
rect 7377 15651 7435 15657
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 8570 15648 8576 15700
rect 8628 15688 8634 15700
rect 8628 15660 8800 15688
rect 8628 15648 8634 15660
rect 4062 15620 4068 15632
rect 3436 15592 4068 15620
rect 4062 15580 4068 15592
rect 4120 15580 4126 15632
rect 5442 15580 5448 15632
rect 5500 15620 5506 15632
rect 5813 15623 5871 15629
rect 5813 15620 5825 15623
rect 5500 15592 5825 15620
rect 5500 15580 5506 15592
rect 5813 15589 5825 15592
rect 5859 15589 5871 15623
rect 5813 15583 5871 15589
rect 3510 15552 3516 15564
rect 2056 15524 3516 15552
rect 2056 15493 2084 15524
rect 1581 15487 1639 15493
rect 1581 15453 1593 15487
rect 1627 15453 1639 15487
rect 1581 15447 1639 15453
rect 2041 15487 2099 15493
rect 2041 15453 2053 15487
rect 2087 15453 2099 15487
rect 2041 15447 2099 15453
rect 1596 15360 1624 15447
rect 2222 15444 2228 15496
rect 2280 15484 2286 15496
rect 2608 15493 2636 15524
rect 3510 15512 3516 15524
rect 3568 15512 3574 15564
rect 4246 15512 4252 15564
rect 4304 15552 4310 15564
rect 8772 15561 8800 15660
rect 11974 15648 11980 15700
rect 12032 15648 12038 15700
rect 13449 15691 13507 15697
rect 13449 15657 13461 15691
rect 13495 15688 13507 15691
rect 13722 15688 13728 15700
rect 13495 15660 13728 15688
rect 13495 15657 13507 15660
rect 13449 15651 13507 15657
rect 13722 15648 13728 15660
rect 13780 15648 13786 15700
rect 14369 15691 14427 15697
rect 14369 15657 14381 15691
rect 14415 15688 14427 15691
rect 15378 15688 15384 15700
rect 14415 15660 15384 15688
rect 14415 15657 14427 15660
rect 14369 15651 14427 15657
rect 15378 15648 15384 15660
rect 15436 15648 15442 15700
rect 15470 15648 15476 15700
rect 15528 15688 15534 15700
rect 15528 15660 16068 15688
rect 15528 15648 15534 15660
rect 16040 15620 16068 15660
rect 16114 15648 16120 15700
rect 16172 15688 16178 15700
rect 17126 15688 17132 15700
rect 16172 15660 17132 15688
rect 16172 15648 16178 15660
rect 17126 15648 17132 15660
rect 17184 15648 17190 15700
rect 19334 15688 19340 15700
rect 17696 15660 19340 15688
rect 17034 15620 17040 15632
rect 16040 15592 17040 15620
rect 17034 15580 17040 15592
rect 17092 15580 17098 15632
rect 4433 15555 4491 15561
rect 4433 15552 4445 15555
rect 4304 15524 4445 15552
rect 4304 15512 4310 15524
rect 4433 15521 4445 15524
rect 4479 15521 4491 15555
rect 4433 15515 4491 15521
rect 8757 15555 8815 15561
rect 8757 15521 8769 15555
rect 8803 15521 8815 15555
rect 8757 15515 8815 15521
rect 10502 15512 10508 15564
rect 10560 15552 10566 15564
rect 10597 15555 10655 15561
rect 10597 15552 10609 15555
rect 10560 15524 10609 15552
rect 10560 15512 10566 15524
rect 10597 15521 10609 15524
rect 10643 15521 10655 15555
rect 14366 15552 14372 15564
rect 10597 15515 10655 15521
rect 13924 15524 14372 15552
rect 2317 15487 2375 15493
rect 2317 15484 2329 15487
rect 2280 15456 2329 15484
rect 2280 15444 2286 15456
rect 2317 15453 2329 15456
rect 2363 15453 2375 15487
rect 2317 15447 2375 15453
rect 2593 15487 2651 15493
rect 2593 15453 2605 15487
rect 2639 15453 2651 15487
rect 2593 15447 2651 15453
rect 2685 15487 2743 15493
rect 2685 15453 2697 15487
rect 2731 15453 2743 15487
rect 2685 15447 2743 15453
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 3602 15484 3608 15496
rect 3099 15456 3608 15484
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 1854 15376 1860 15428
rect 1912 15416 1918 15428
rect 2501 15419 2559 15425
rect 2501 15416 2513 15419
rect 1912 15388 2513 15416
rect 1912 15376 1918 15388
rect 2501 15385 2513 15388
rect 2547 15385 2559 15419
rect 2501 15379 2559 15385
rect 1578 15308 1584 15360
rect 1636 15308 1642 15360
rect 1762 15308 1768 15360
rect 1820 15348 1826 15360
rect 1949 15351 2007 15357
rect 1949 15348 1961 15351
rect 1820 15320 1961 15348
rect 1820 15308 1826 15320
rect 1949 15317 1961 15320
rect 1995 15317 2007 15351
rect 1949 15311 2007 15317
rect 2130 15308 2136 15360
rect 2188 15308 2194 15360
rect 2406 15308 2412 15360
rect 2464 15348 2470 15360
rect 2700 15348 2728 15447
rect 3602 15444 3608 15456
rect 3660 15444 3666 15496
rect 3694 15444 3700 15496
rect 3752 15444 3758 15496
rect 3970 15444 3976 15496
rect 4028 15484 4034 15496
rect 4065 15487 4123 15493
rect 4065 15484 4077 15487
rect 4028 15456 4077 15484
rect 4028 15444 4034 15456
rect 4065 15453 4077 15456
rect 4111 15453 4123 15487
rect 4065 15447 4123 15453
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15484 4215 15487
rect 4522 15484 4528 15496
rect 4203 15456 4528 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 4522 15444 4528 15456
rect 4580 15444 4586 15496
rect 5905 15487 5963 15493
rect 5905 15484 5917 15487
rect 4632 15456 5917 15484
rect 2464 15320 2728 15348
rect 2777 15351 2835 15357
rect 2464 15308 2470 15320
rect 2777 15317 2789 15351
rect 2823 15348 2835 15351
rect 3326 15348 3332 15360
rect 2823 15320 3332 15348
rect 2823 15317 2835 15320
rect 2777 15311 2835 15317
rect 3326 15308 3332 15320
rect 3384 15308 3390 15360
rect 3712 15348 3740 15444
rect 4249 15419 4307 15425
rect 4249 15385 4261 15419
rect 4295 15416 4307 15419
rect 4632 15416 4660 15456
rect 5905 15453 5917 15456
rect 5951 15453 5963 15487
rect 5905 15447 5963 15453
rect 9858 15444 9864 15496
rect 9916 15484 9922 15496
rect 10870 15493 10876 15496
rect 10413 15487 10471 15493
rect 10413 15484 10425 15487
rect 9916 15456 10425 15484
rect 9916 15444 9922 15456
rect 10413 15453 10425 15456
rect 10459 15453 10471 15487
rect 10864 15484 10876 15493
rect 10831 15456 10876 15484
rect 10413 15447 10471 15453
rect 10864 15447 10876 15456
rect 10870 15444 10876 15447
rect 10928 15444 10934 15496
rect 12066 15444 12072 15496
rect 12124 15444 12130 15496
rect 13924 15493 13952 15524
rect 14366 15512 14372 15524
rect 14424 15512 14430 15564
rect 16482 15552 16488 15564
rect 15672 15524 16488 15552
rect 13909 15487 13967 15493
rect 13909 15453 13921 15487
rect 13955 15453 13967 15487
rect 13909 15447 13967 15453
rect 14277 15487 14335 15493
rect 14277 15453 14289 15487
rect 14323 15484 14335 15487
rect 15672 15484 15700 15524
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 16942 15512 16948 15564
rect 17000 15512 17006 15564
rect 17696 15561 17724 15660
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 18874 15580 18880 15632
rect 18932 15620 18938 15632
rect 20533 15623 20591 15629
rect 20533 15620 20545 15623
rect 18932 15592 20545 15620
rect 18932 15580 18938 15592
rect 20533 15589 20545 15592
rect 20579 15620 20591 15623
rect 21082 15620 21088 15632
rect 20579 15592 21088 15620
rect 20579 15589 20591 15592
rect 20533 15583 20591 15589
rect 21082 15580 21088 15592
rect 21140 15580 21146 15632
rect 17681 15555 17739 15561
rect 17681 15521 17693 15555
rect 17727 15521 17739 15555
rect 17681 15515 17739 15521
rect 22465 15555 22523 15561
rect 22465 15521 22477 15555
rect 22511 15552 22523 15555
rect 23385 15555 23443 15561
rect 23385 15552 23397 15555
rect 22511 15524 23397 15552
rect 22511 15521 22523 15524
rect 22465 15515 22523 15521
rect 23385 15521 23397 15524
rect 23431 15521 23443 15555
rect 23385 15515 23443 15521
rect 14323 15456 15700 15484
rect 15749 15487 15807 15493
rect 14323 15453 14335 15456
rect 14277 15447 14335 15453
rect 15749 15453 15761 15487
rect 15795 15484 15807 15487
rect 16960 15484 16988 15512
rect 15795 15456 16988 15484
rect 15795 15453 15807 15456
rect 15749 15447 15807 15453
rect 17586 15444 17592 15496
rect 17644 15484 17650 15496
rect 19245 15487 19303 15493
rect 19245 15484 19257 15487
rect 17644 15456 19257 15484
rect 17644 15444 17650 15456
rect 19245 15453 19257 15456
rect 19291 15453 19303 15487
rect 19245 15447 19303 15453
rect 22209 15487 22267 15493
rect 22209 15453 22221 15487
rect 22255 15484 22267 15487
rect 22554 15484 22560 15496
rect 22255 15456 22560 15484
rect 22255 15453 22267 15456
rect 22209 15447 22267 15453
rect 22554 15444 22560 15456
rect 22612 15444 22618 15496
rect 22646 15444 22652 15496
rect 22704 15484 22710 15496
rect 23109 15487 23167 15493
rect 23109 15484 23121 15487
rect 22704 15456 23121 15484
rect 22704 15444 22710 15456
rect 23109 15453 23121 15456
rect 23155 15453 23167 15487
rect 23109 15447 23167 15453
rect 23293 15487 23351 15493
rect 23293 15453 23305 15487
rect 23339 15453 23351 15487
rect 23293 15447 23351 15453
rect 4706 15425 4712 15428
rect 4295 15388 4660 15416
rect 4295 15385 4307 15388
rect 4249 15379 4307 15385
rect 4700 15379 4712 15425
rect 4706 15376 4712 15379
rect 4764 15376 4770 15428
rect 6150 15419 6208 15425
rect 6150 15416 6162 15419
rect 4816 15388 6162 15416
rect 4816 15348 4844 15388
rect 6150 15385 6162 15388
rect 6196 15385 6208 15419
rect 6150 15379 6208 15385
rect 8386 15376 8392 15428
rect 8444 15416 8450 15428
rect 8490 15419 8548 15425
rect 8490 15416 8502 15419
rect 8444 15388 8502 15416
rect 8444 15376 8450 15388
rect 8490 15385 8502 15388
rect 8536 15385 8548 15419
rect 8490 15379 8548 15385
rect 9950 15376 9956 15428
rect 10008 15416 10014 15428
rect 12342 15425 12348 15428
rect 10146 15419 10204 15425
rect 10146 15416 10158 15419
rect 10008 15388 10158 15416
rect 10008 15376 10014 15388
rect 10146 15385 10158 15388
rect 10192 15385 10204 15419
rect 10146 15379 10204 15385
rect 12336 15379 12348 15425
rect 12342 15376 12348 15379
rect 12400 15376 12406 15428
rect 14185 15419 14243 15425
rect 14185 15385 14197 15419
rect 14231 15416 14243 15419
rect 15194 15416 15200 15428
rect 14231 15388 15200 15416
rect 14231 15385 14243 15388
rect 14185 15379 14243 15385
rect 15194 15376 15200 15388
rect 15252 15376 15258 15428
rect 15470 15376 15476 15428
rect 15528 15425 15534 15428
rect 15528 15419 15562 15425
rect 15550 15385 15562 15419
rect 15841 15419 15899 15425
rect 15841 15416 15853 15419
rect 15528 15379 15562 15385
rect 15672 15388 15853 15416
rect 15528 15376 15534 15379
rect 3712 15320 4844 15348
rect 9033 15351 9091 15357
rect 9033 15317 9045 15351
rect 9079 15348 9091 15351
rect 9214 15348 9220 15360
rect 9079 15320 9220 15348
rect 9079 15317 9091 15320
rect 9033 15311 9091 15317
rect 9214 15308 9220 15320
rect 9272 15308 9278 15360
rect 13814 15308 13820 15360
rect 13872 15308 13878 15360
rect 14550 15308 14556 15360
rect 14608 15348 14614 15360
rect 15672 15348 15700 15388
rect 15841 15385 15853 15388
rect 15887 15385 15899 15419
rect 15841 15379 15899 15385
rect 17948 15419 18006 15425
rect 17948 15385 17960 15419
rect 17994 15416 18006 15419
rect 18138 15416 18144 15428
rect 17994 15388 18144 15416
rect 17994 15385 18006 15388
rect 17948 15379 18006 15385
rect 18138 15376 18144 15388
rect 18196 15376 18202 15428
rect 19518 15376 19524 15428
rect 19576 15416 19582 15428
rect 23014 15416 23020 15428
rect 19576 15388 23020 15416
rect 19576 15376 19582 15388
rect 23014 15376 23020 15388
rect 23072 15376 23078 15428
rect 23308 15416 23336 15447
rect 23124 15388 23336 15416
rect 23124 15360 23152 15388
rect 14608 15320 15700 15348
rect 19061 15351 19119 15357
rect 14608 15308 14614 15320
rect 19061 15317 19073 15351
rect 19107 15348 19119 15351
rect 19610 15348 19616 15360
rect 19107 15320 19616 15348
rect 19107 15317 19119 15320
rect 19061 15311 19119 15317
rect 19610 15308 19616 15320
rect 19668 15308 19674 15360
rect 21085 15351 21143 15357
rect 21085 15317 21097 15351
rect 21131 15348 21143 15351
rect 21358 15348 21364 15360
rect 21131 15320 21364 15348
rect 21131 15317 21143 15320
rect 21085 15311 21143 15317
rect 21358 15308 21364 15320
rect 21416 15308 21422 15360
rect 22554 15308 22560 15360
rect 22612 15308 22618 15360
rect 23106 15308 23112 15360
rect 23164 15308 23170 15360
rect 1104 15258 23828 15280
rect 1104 15206 2658 15258
rect 2710 15206 2722 15258
rect 2774 15206 2786 15258
rect 2838 15206 2850 15258
rect 2902 15206 2914 15258
rect 2966 15206 2978 15258
rect 3030 15206 8658 15258
rect 8710 15206 8722 15258
rect 8774 15206 8786 15258
rect 8838 15206 8850 15258
rect 8902 15206 8914 15258
rect 8966 15206 8978 15258
rect 9030 15206 14658 15258
rect 14710 15206 14722 15258
rect 14774 15206 14786 15258
rect 14838 15206 14850 15258
rect 14902 15206 14914 15258
rect 14966 15206 14978 15258
rect 15030 15206 20658 15258
rect 20710 15206 20722 15258
rect 20774 15206 20786 15258
rect 20838 15206 20850 15258
rect 20902 15206 20914 15258
rect 20966 15206 20978 15258
rect 21030 15206 23828 15258
rect 1104 15184 23828 15206
rect 1578 15104 1584 15156
rect 1636 15144 1642 15156
rect 3234 15144 3240 15156
rect 1636 15116 3240 15144
rect 1636 15104 1642 15116
rect 3234 15104 3240 15116
rect 3292 15104 3298 15156
rect 4430 15144 4436 15156
rect 3344 15116 4436 15144
rect 1596 15017 1624 15104
rect 2124 15079 2182 15085
rect 2124 15045 2136 15079
rect 2170 15076 2182 15079
rect 3050 15076 3056 15088
rect 2170 15048 3056 15076
rect 2170 15045 2182 15048
rect 2124 15039 2182 15045
rect 3050 15036 3056 15048
rect 3108 15036 3114 15088
rect 1581 15011 1639 15017
rect 1581 14977 1593 15011
rect 1627 14977 1639 15011
rect 1581 14971 1639 14977
rect 3142 14968 3148 15020
rect 3200 15008 3206 15020
rect 3344 15017 3372 15116
rect 4430 15104 4436 15116
rect 4488 15104 4494 15156
rect 5074 15144 5080 15156
rect 4540 15116 5080 15144
rect 3694 15036 3700 15088
rect 3752 15076 3758 15088
rect 4540 15076 4568 15116
rect 5074 15104 5080 15116
rect 5132 15104 5138 15156
rect 6086 15104 6092 15156
rect 6144 15144 6150 15156
rect 6181 15147 6239 15153
rect 6181 15144 6193 15147
rect 6144 15116 6193 15144
rect 6144 15104 6150 15116
rect 6181 15113 6193 15116
rect 6227 15113 6239 15147
rect 6181 15107 6239 15113
rect 7098 15104 7104 15156
rect 7156 15144 7162 15156
rect 7745 15147 7803 15153
rect 7745 15144 7757 15147
rect 7156 15116 7757 15144
rect 7156 15104 7162 15116
rect 7745 15113 7757 15116
rect 7791 15113 7803 15147
rect 7745 15107 7803 15113
rect 8297 15147 8355 15153
rect 8297 15113 8309 15147
rect 8343 15144 8355 15147
rect 8478 15144 8484 15156
rect 8343 15116 8484 15144
rect 8343 15113 8355 15116
rect 8297 15107 8355 15113
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 9769 15147 9827 15153
rect 9769 15113 9781 15147
rect 9815 15144 9827 15147
rect 12066 15144 12072 15156
rect 9815 15116 12072 15144
rect 9815 15113 9827 15116
rect 9769 15107 9827 15113
rect 12066 15104 12072 15116
rect 12124 15104 12130 15156
rect 12345 15147 12403 15153
rect 12345 15113 12357 15147
rect 12391 15113 12403 15147
rect 12345 15107 12403 15113
rect 3752 15048 4568 15076
rect 3752 15036 3758 15048
rect 4614 15036 4620 15088
rect 4672 15076 4678 15088
rect 11054 15076 11060 15088
rect 4672 15048 6408 15076
rect 4672 15036 4678 15048
rect 3329 15011 3387 15017
rect 3329 15008 3341 15011
rect 3200 14980 3341 15008
rect 3200 14968 3206 14980
rect 3329 14977 3341 14980
rect 3375 14977 3387 15011
rect 3585 15011 3643 15017
rect 3585 15008 3597 15011
rect 3329 14971 3387 14977
rect 3436 14980 3597 15008
rect 1854 14900 1860 14952
rect 1912 14900 1918 14952
rect 3436 14940 3464 14980
rect 3585 14977 3597 14980
rect 3631 14977 3643 15011
rect 3585 14971 3643 14977
rect 4154 14968 4160 15020
rect 4212 15008 4218 15020
rect 6380 15017 6408 15048
rect 9692 15048 11060 15076
rect 4801 15011 4859 15017
rect 4801 15008 4813 15011
rect 4212 14980 4813 15008
rect 4212 14968 4218 14980
rect 4801 14977 4813 14980
rect 4847 14977 4859 15011
rect 5057 15011 5115 15017
rect 5057 15008 5069 15011
rect 4801 14971 4859 14977
rect 4908 14980 5069 15008
rect 4908 14940 4936 14980
rect 5057 14977 5069 14980
rect 5103 14977 5115 15011
rect 5057 14971 5115 14977
rect 6365 15011 6423 15017
rect 6365 14977 6377 15011
rect 6411 14977 6423 15011
rect 6621 15011 6679 15017
rect 6621 15008 6633 15011
rect 6365 14971 6423 14977
rect 6472 14980 6633 15008
rect 6472 14940 6500 14980
rect 6621 14977 6633 14980
rect 6667 14977 6679 15011
rect 6621 14971 6679 14977
rect 9582 14968 9588 15020
rect 9640 14968 9646 15020
rect 9692 15017 9720 15048
rect 11054 15036 11060 15048
rect 11112 15036 11118 15088
rect 9677 15011 9735 15017
rect 9677 14977 9689 15011
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 9766 14968 9772 15020
rect 9824 15008 9830 15020
rect 9953 15011 10011 15017
rect 9953 15008 9965 15011
rect 9824 14980 9965 15008
rect 9824 14968 9830 14980
rect 9953 14977 9965 14980
rect 9999 14977 10011 15011
rect 9953 14971 10011 14977
rect 10220 15011 10278 15017
rect 10220 14977 10232 15011
rect 10266 15008 10278 15011
rect 10778 15008 10784 15020
rect 10266 14980 10784 15008
rect 10266 14977 10278 14980
rect 10220 14971 10278 14977
rect 10778 14968 10784 14980
rect 10836 14968 10842 15020
rect 12253 15011 12311 15017
rect 12253 14977 12265 15011
rect 12299 15008 12311 15011
rect 12360 15008 12388 15107
rect 14366 15104 14372 15156
rect 14424 15144 14430 15156
rect 14424 15116 20024 15144
rect 14424 15104 14430 15116
rect 13446 15036 13452 15088
rect 13504 15085 13510 15088
rect 13504 15079 13538 15085
rect 13526 15045 13538 15079
rect 13504 15039 13538 15045
rect 15657 15079 15715 15085
rect 15657 15045 15669 15079
rect 15703 15076 15715 15079
rect 17586 15076 17592 15088
rect 15703 15048 17592 15076
rect 15703 15045 15715 15048
rect 15657 15039 15715 15045
rect 13504 15036 13510 15039
rect 17586 15036 17592 15048
rect 17644 15036 17650 15088
rect 19242 15076 19248 15088
rect 17696 15048 19248 15076
rect 17696 15020 17724 15048
rect 19242 15036 19248 15048
rect 19300 15036 19306 15088
rect 19702 15036 19708 15088
rect 19760 15076 19766 15088
rect 19858 15079 19916 15085
rect 19858 15076 19870 15079
rect 19760 15048 19870 15076
rect 19760 15036 19766 15048
rect 19858 15045 19870 15048
rect 19904 15045 19916 15079
rect 19858 15039 19916 15045
rect 12299 14980 12388 15008
rect 13725 15011 13783 15017
rect 12299 14977 12311 14980
rect 12253 14971 12311 14977
rect 13725 14977 13737 15011
rect 13771 15008 13783 15011
rect 13814 15008 13820 15020
rect 13771 14980 13820 15008
rect 13771 14977 13783 14980
rect 13725 14971 13783 14977
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 16574 14968 16580 15020
rect 16632 15008 16638 15020
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 16632 14980 16681 15008
rect 16632 14968 16638 14980
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 16936 15011 16994 15017
rect 16936 14977 16948 15011
rect 16982 15008 16994 15011
rect 17218 15008 17224 15020
rect 16982 14980 17224 15008
rect 16982 14977 16994 14980
rect 16936 14971 16994 14977
rect 17218 14968 17224 14980
rect 17276 14968 17282 15020
rect 17678 14968 17684 15020
rect 17736 14968 17742 15020
rect 17954 14968 17960 15020
rect 18012 15008 18018 15020
rect 18141 15011 18199 15017
rect 18141 15008 18153 15011
rect 18012 14980 18153 15008
rect 18012 14968 18018 14980
rect 18141 14977 18153 14980
rect 18187 14977 18199 15011
rect 18397 15011 18455 15017
rect 18397 15008 18409 15011
rect 18141 14971 18199 14977
rect 18248 14980 18409 15008
rect 3252 14912 3464 14940
rect 4724 14912 4936 14940
rect 5828 14912 6500 14940
rect 3252 14881 3280 14912
rect 4724 14881 4752 14912
rect 3237 14875 3295 14881
rect 3237 14841 3249 14875
rect 3283 14841 3295 14875
rect 3237 14835 3295 14841
rect 4709 14875 4767 14881
rect 4709 14841 4721 14875
rect 4755 14841 4767 14875
rect 4709 14835 4767 14841
rect 1670 14764 1676 14816
rect 1728 14764 1734 14816
rect 2130 14764 2136 14816
rect 2188 14804 2194 14816
rect 2590 14804 2596 14816
rect 2188 14776 2596 14804
rect 2188 14764 2194 14776
rect 2590 14764 2596 14776
rect 2648 14764 2654 14816
rect 3602 14764 3608 14816
rect 3660 14804 3666 14816
rect 5828 14804 5856 14912
rect 16298 14900 16304 14952
rect 16356 14900 16362 14952
rect 18248 14940 18276 14980
rect 18397 14977 18409 14980
rect 18443 14977 18455 15011
rect 18397 14971 18455 14977
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 19613 15011 19671 15017
rect 19613 15008 19625 15011
rect 19484 14980 19625 15008
rect 19484 14968 19490 14980
rect 19613 14977 19625 14980
rect 19659 14977 19671 15011
rect 19996 15008 20024 15116
rect 21082 15104 21088 15156
rect 21140 15104 21146 15156
rect 21821 15147 21879 15153
rect 21821 15113 21833 15147
rect 21867 15144 21879 15147
rect 22094 15144 22100 15156
rect 21867 15116 22100 15144
rect 21867 15113 21879 15116
rect 21821 15107 21879 15113
rect 22094 15104 22100 15116
rect 22152 15104 22158 15156
rect 21100 15076 21128 15104
rect 21100 15048 21588 15076
rect 21560 15017 21588 15048
rect 21634 15036 21640 15088
rect 21692 15076 21698 15088
rect 21692 15048 23336 15076
rect 21692 15036 21698 15048
rect 23308 15020 23336 15048
rect 21085 15011 21143 15017
rect 21085 15008 21097 15011
rect 19996 14980 21097 15008
rect 19613 14971 19671 14977
rect 21085 14977 21097 14980
rect 21131 14977 21143 15011
rect 21085 14971 21143 14977
rect 21545 15011 21603 15017
rect 21545 14977 21557 15011
rect 21591 14977 21603 15011
rect 22370 15008 22376 15020
rect 21545 14971 21603 14977
rect 22066 14980 22376 15008
rect 17696 14912 18276 14940
rect 10980 14844 12434 14872
rect 10980 14816 11008 14844
rect 3660 14776 5856 14804
rect 3660 14764 3666 14776
rect 6362 14764 6368 14816
rect 6420 14804 6426 14816
rect 9950 14804 9956 14816
rect 6420 14776 9956 14804
rect 6420 14764 6426 14776
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 10962 14764 10968 14816
rect 11020 14764 11026 14816
rect 11330 14764 11336 14816
rect 11388 14764 11394 14816
rect 11606 14764 11612 14816
rect 11664 14764 11670 14816
rect 12406 14804 12434 14844
rect 14366 14804 14372 14816
rect 12406 14776 14372 14804
rect 14366 14764 14372 14776
rect 14424 14764 14430 14816
rect 15746 14764 15752 14816
rect 15804 14764 15810 14816
rect 16482 14764 16488 14816
rect 16540 14804 16546 14816
rect 17696 14804 17724 14912
rect 19518 14900 19524 14952
rect 19576 14900 19582 14952
rect 20622 14900 20628 14952
rect 20680 14940 20686 14952
rect 22066 14940 22094 14980
rect 22370 14968 22376 14980
rect 22428 14968 22434 15020
rect 22945 15011 23003 15017
rect 22945 14977 22957 15011
rect 22991 15008 23003 15011
rect 22991 14980 23152 15008
rect 22991 14977 23003 14980
rect 22945 14971 23003 14977
rect 20680 14912 22094 14940
rect 23124 14940 23152 14980
rect 23198 14968 23204 15020
rect 23256 14968 23262 15020
rect 23290 14968 23296 15020
rect 23348 14968 23354 15020
rect 23124 14912 23244 14940
rect 20680 14900 20686 14912
rect 19536 14872 19564 14900
rect 23216 14884 23244 14912
rect 19444 14844 19564 14872
rect 20993 14875 21051 14881
rect 16540 14776 17724 14804
rect 18049 14807 18107 14813
rect 16540 14764 16546 14776
rect 18049 14773 18061 14807
rect 18095 14804 18107 14807
rect 19444 14804 19472 14844
rect 20993 14841 21005 14875
rect 21039 14872 21051 14875
rect 21039 14844 22094 14872
rect 21039 14841 21051 14844
rect 20993 14835 21051 14841
rect 18095 14776 19472 14804
rect 19521 14807 19579 14813
rect 18095 14773 18107 14776
rect 18049 14767 18107 14773
rect 19521 14773 19533 14807
rect 19567 14804 19579 14807
rect 19794 14804 19800 14816
rect 19567 14776 19800 14804
rect 19567 14773 19579 14776
rect 19521 14767 19579 14773
rect 19794 14764 19800 14776
rect 19852 14764 19858 14816
rect 20530 14764 20536 14816
rect 20588 14804 20594 14816
rect 21177 14807 21235 14813
rect 21177 14804 21189 14807
rect 20588 14776 21189 14804
rect 20588 14764 20594 14776
rect 21177 14773 21189 14776
rect 21223 14773 21235 14807
rect 21177 14767 21235 14773
rect 21266 14764 21272 14816
rect 21324 14804 21330 14816
rect 21453 14807 21511 14813
rect 21453 14804 21465 14807
rect 21324 14776 21465 14804
rect 21324 14764 21330 14776
rect 21453 14773 21465 14776
rect 21499 14773 21511 14807
rect 22066 14804 22094 14844
rect 23198 14832 23204 14884
rect 23256 14832 23262 14884
rect 22278 14804 22284 14816
rect 22066 14776 22284 14804
rect 21453 14767 21511 14773
rect 22278 14764 22284 14776
rect 22336 14764 22342 14816
rect 22462 14764 22468 14816
rect 22520 14804 22526 14816
rect 23385 14807 23443 14813
rect 23385 14804 23397 14807
rect 22520 14776 23397 14804
rect 22520 14764 22526 14776
rect 23385 14773 23397 14776
rect 23431 14773 23443 14807
rect 23385 14767 23443 14773
rect 1104 14714 23828 14736
rect 1104 14662 1918 14714
rect 1970 14662 1982 14714
rect 2034 14662 2046 14714
rect 2098 14662 2110 14714
rect 2162 14662 2174 14714
rect 2226 14662 2238 14714
rect 2290 14662 7918 14714
rect 7970 14662 7982 14714
rect 8034 14662 8046 14714
rect 8098 14662 8110 14714
rect 8162 14662 8174 14714
rect 8226 14662 8238 14714
rect 8290 14662 13918 14714
rect 13970 14662 13982 14714
rect 14034 14662 14046 14714
rect 14098 14662 14110 14714
rect 14162 14662 14174 14714
rect 14226 14662 14238 14714
rect 14290 14662 19918 14714
rect 19970 14662 19982 14714
rect 20034 14662 20046 14714
rect 20098 14662 20110 14714
rect 20162 14662 20174 14714
rect 20226 14662 20238 14714
rect 20290 14662 23828 14714
rect 1104 14640 23828 14662
rect 1670 14560 1676 14612
rect 1728 14600 1734 14612
rect 1728 14572 6776 14600
rect 1728 14560 1734 14572
rect 3510 14532 3516 14544
rect 2746 14504 3516 14532
rect 2317 14467 2375 14473
rect 2317 14433 2329 14467
rect 2363 14464 2375 14467
rect 2746 14464 2774 14504
rect 3510 14492 3516 14504
rect 3568 14492 3574 14544
rect 3602 14492 3608 14544
rect 3660 14492 3666 14544
rect 5074 14492 5080 14544
rect 5132 14532 5138 14544
rect 5261 14535 5319 14541
rect 5261 14532 5273 14535
rect 5132 14504 5273 14532
rect 5132 14492 5138 14504
rect 5261 14501 5273 14504
rect 5307 14501 5319 14535
rect 5261 14495 5319 14501
rect 5353 14535 5411 14541
rect 5353 14501 5365 14535
rect 5399 14501 5411 14535
rect 5353 14495 5411 14501
rect 2363 14436 2774 14464
rect 2363 14433 2375 14436
rect 2317 14427 2375 14433
rect 3326 14424 3332 14476
rect 3384 14464 3390 14476
rect 3881 14467 3939 14473
rect 3881 14464 3893 14467
rect 3384 14436 3893 14464
rect 3384 14424 3390 14436
rect 3881 14433 3893 14436
rect 3927 14433 3939 14467
rect 3881 14427 3939 14433
rect 2041 14399 2099 14405
rect 2041 14365 2053 14399
rect 2087 14396 2099 14399
rect 3053 14399 3111 14405
rect 2087 14368 2774 14396
rect 2087 14365 2099 14368
rect 2041 14359 2099 14365
rect 1302 14288 1308 14340
rect 1360 14328 1366 14340
rect 1489 14331 1547 14337
rect 1489 14328 1501 14331
rect 1360 14300 1501 14328
rect 1360 14288 1366 14300
rect 1489 14297 1501 14300
rect 1535 14297 1547 14331
rect 1489 14291 1547 14297
rect 2130 14288 2136 14340
rect 2188 14328 2194 14340
rect 2590 14328 2596 14340
rect 2188 14300 2596 14328
rect 2188 14288 2194 14300
rect 2590 14288 2596 14300
rect 2648 14288 2654 14340
rect 2746 14260 2774 14368
rect 3053 14365 3065 14399
rect 3099 14396 3111 14399
rect 5368 14396 5396 14495
rect 6748 14473 6776 14572
rect 9674 14560 9680 14612
rect 9732 14560 9738 14612
rect 11974 14560 11980 14612
rect 12032 14600 12038 14612
rect 16298 14600 16304 14612
rect 12032 14572 16304 14600
rect 12032 14560 12038 14572
rect 16298 14560 16304 14572
rect 16356 14560 16362 14612
rect 17034 14560 17040 14612
rect 17092 14560 17098 14612
rect 20530 14600 20536 14612
rect 18432 14572 20536 14600
rect 6733 14467 6791 14473
rect 6733 14433 6745 14467
rect 6779 14433 6791 14467
rect 6733 14427 6791 14433
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14464 9643 14467
rect 9692 14464 9720 14560
rect 13814 14532 13820 14544
rect 9631 14436 9720 14464
rect 13004 14504 13820 14532
rect 9631 14433 9643 14436
rect 9585 14427 9643 14433
rect 3099 14368 5396 14396
rect 3099 14365 3111 14368
rect 3053 14359 3111 14365
rect 6454 14356 6460 14408
rect 6512 14405 6518 14408
rect 6512 14396 6524 14405
rect 9677 14399 9735 14405
rect 6512 14368 6557 14396
rect 6512 14359 6524 14368
rect 9677 14365 9689 14399
rect 9723 14396 9735 14399
rect 9766 14396 9772 14408
rect 9723 14368 9772 14396
rect 9723 14365 9735 14368
rect 9677 14359 9735 14365
rect 6512 14356 6518 14359
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 13004 14396 13032 14504
rect 13814 14492 13820 14504
rect 13872 14492 13878 14544
rect 13081 14467 13139 14473
rect 13081 14433 13093 14467
rect 13127 14464 13139 14467
rect 14093 14467 14151 14473
rect 14093 14464 14105 14467
rect 13127 14436 14105 14464
rect 13127 14433 13139 14436
rect 13081 14427 13139 14433
rect 14093 14433 14105 14436
rect 14139 14433 14151 14467
rect 14093 14427 14151 14433
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 18432 14473 18460 14572
rect 20530 14560 20536 14572
rect 20588 14560 20594 14612
rect 22646 14600 22652 14612
rect 21192 14572 22652 14600
rect 18877 14535 18935 14541
rect 18877 14501 18889 14535
rect 18923 14532 18935 14535
rect 20625 14535 20683 14541
rect 18923 14504 19196 14532
rect 18923 14501 18935 14504
rect 18877 14495 18935 14501
rect 15565 14467 15623 14473
rect 15565 14464 15577 14467
rect 15252 14436 15577 14464
rect 15252 14424 15258 14436
rect 15565 14433 15577 14436
rect 15611 14433 15623 14467
rect 15565 14427 15623 14433
rect 18417 14467 18475 14473
rect 18417 14433 18429 14467
rect 18463 14433 18475 14467
rect 18417 14427 18475 14433
rect 18509 14467 18567 14473
rect 18509 14433 18521 14467
rect 18555 14464 18567 14467
rect 18598 14464 18604 14476
rect 18555 14436 18604 14464
rect 18555 14433 18567 14436
rect 18509 14427 18567 14433
rect 18598 14424 18604 14436
rect 18656 14424 18662 14476
rect 13173 14399 13231 14405
rect 13173 14396 13185 14399
rect 13004 14368 13185 14396
rect 13173 14365 13185 14368
rect 13219 14365 13231 14399
rect 13173 14359 13231 14365
rect 13354 14356 13360 14408
rect 13412 14356 13418 14408
rect 13909 14399 13967 14405
rect 13909 14365 13921 14399
rect 13955 14396 13967 14399
rect 14349 14399 14407 14405
rect 14349 14396 14361 14399
rect 13955 14368 14361 14396
rect 13955 14365 13967 14368
rect 13909 14359 13967 14365
rect 14349 14365 14361 14368
rect 14395 14365 14407 14399
rect 14349 14359 14407 14365
rect 15378 14356 15384 14408
rect 15436 14396 15442 14408
rect 15821 14399 15879 14405
rect 15821 14396 15833 14399
rect 15436 14368 15833 14396
rect 15436 14356 15442 14368
rect 15821 14365 15833 14368
rect 15867 14365 15879 14399
rect 15821 14359 15879 14365
rect 17126 14356 17132 14408
rect 17184 14396 17190 14408
rect 18150 14399 18208 14405
rect 18150 14396 18162 14399
rect 17184 14368 18162 14396
rect 17184 14356 17190 14368
rect 18150 14365 18162 14368
rect 18196 14365 18208 14399
rect 18150 14359 18208 14365
rect 18432 14368 19104 14396
rect 2869 14331 2927 14337
rect 2869 14297 2881 14331
rect 2915 14328 2927 14331
rect 3418 14328 3424 14340
rect 2915 14300 3424 14328
rect 2915 14297 2927 14300
rect 2869 14291 2927 14297
rect 3418 14288 3424 14300
rect 3476 14288 3482 14340
rect 3878 14328 3884 14340
rect 3620 14300 3884 14328
rect 3620 14260 3648 14300
rect 3878 14288 3884 14300
rect 3936 14288 3942 14340
rect 4148 14331 4206 14337
rect 4148 14297 4160 14331
rect 4194 14328 4206 14331
rect 4430 14328 4436 14340
rect 4194 14300 4436 14328
rect 4194 14297 4206 14300
rect 4148 14291 4206 14297
rect 4430 14288 4436 14300
rect 4488 14288 4494 14340
rect 4706 14288 4712 14340
rect 4764 14288 4770 14340
rect 9950 14337 9956 14340
rect 8573 14331 8631 14337
rect 8573 14297 8585 14331
rect 8619 14328 8631 14331
rect 8619 14300 9536 14328
rect 8619 14297 8631 14300
rect 8573 14291 8631 14297
rect 2746 14232 3648 14260
rect 3694 14220 3700 14272
rect 3752 14260 3758 14272
rect 4724 14260 4752 14288
rect 9508 14272 9536 14300
rect 9944 14291 9956 14337
rect 9950 14288 9956 14291
rect 10008 14288 10014 14340
rect 12158 14328 12164 14340
rect 11072 14300 12164 14328
rect 3752 14232 4752 14260
rect 3752 14220 3758 14232
rect 7098 14220 7104 14272
rect 7156 14220 7162 14272
rect 7282 14220 7288 14272
rect 7340 14260 7346 14272
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 7340 14232 8953 14260
rect 7340 14220 7346 14232
rect 8941 14229 8953 14232
rect 8987 14229 8999 14263
rect 8941 14223 8999 14229
rect 9490 14220 9496 14272
rect 9548 14220 9554 14272
rect 11072 14269 11100 14300
rect 12158 14288 12164 14300
rect 12216 14288 12222 14340
rect 12897 14331 12955 14337
rect 12897 14297 12909 14331
rect 12943 14328 12955 14331
rect 14182 14328 14188 14340
rect 12943 14300 14188 14328
rect 12943 14297 12955 14300
rect 12897 14291 12955 14297
rect 14182 14288 14188 14300
rect 14240 14288 14246 14340
rect 18432 14328 18460 14368
rect 15488 14300 18460 14328
rect 11057 14263 11115 14269
rect 11057 14229 11069 14263
rect 11103 14229 11115 14263
rect 11057 14223 11115 14229
rect 11146 14220 11152 14272
rect 11204 14260 11210 14272
rect 11425 14263 11483 14269
rect 11425 14260 11437 14263
rect 11204 14232 11437 14260
rect 11204 14220 11210 14232
rect 11425 14229 11437 14232
rect 11471 14260 11483 14263
rect 13538 14260 13544 14272
rect 11471 14232 13544 14260
rect 11471 14229 11483 14232
rect 11425 14223 11483 14229
rect 13538 14220 13544 14232
rect 13596 14220 13602 14272
rect 15488 14269 15516 14300
rect 15473 14263 15531 14269
rect 15473 14229 15485 14263
rect 15519 14229 15531 14263
rect 15473 14223 15531 14229
rect 16390 14220 16396 14272
rect 16448 14260 16454 14272
rect 16945 14263 17003 14269
rect 16945 14260 16957 14263
rect 16448 14232 16957 14260
rect 16448 14220 16454 14232
rect 16945 14229 16957 14232
rect 16991 14229 17003 14263
rect 16945 14223 17003 14229
rect 18046 14220 18052 14272
rect 18104 14260 18110 14272
rect 18598 14260 18604 14272
rect 18104 14232 18604 14260
rect 18104 14220 18110 14232
rect 18598 14220 18604 14232
rect 18656 14220 18662 14272
rect 18966 14220 18972 14272
rect 19024 14220 19030 14272
rect 19076 14260 19104 14368
rect 19168 14328 19196 14504
rect 20625 14501 20637 14535
rect 20671 14532 20683 14535
rect 21192 14532 21220 14572
rect 22646 14560 22652 14572
rect 22704 14560 22710 14612
rect 20671 14504 21220 14532
rect 20671 14501 20683 14504
rect 20625 14495 20683 14501
rect 22020 14436 23060 14464
rect 19245 14399 19303 14405
rect 19245 14365 19257 14399
rect 19291 14396 19303 14399
rect 20438 14396 20444 14408
rect 19291 14368 20444 14396
rect 19291 14365 19303 14368
rect 19245 14359 19303 14365
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 22020 14396 22048 14436
rect 20732 14368 22048 14396
rect 19334 14328 19340 14340
rect 19168 14300 19340 14328
rect 19334 14288 19340 14300
rect 19392 14288 19398 14340
rect 19512 14331 19570 14337
rect 19512 14297 19524 14331
rect 19558 14328 19570 14331
rect 19794 14328 19800 14340
rect 19558 14300 19800 14328
rect 19558 14297 19570 14300
rect 19512 14291 19570 14297
rect 19794 14288 19800 14300
rect 19852 14288 19858 14340
rect 20622 14260 20628 14272
rect 19076 14232 20628 14260
rect 20622 14220 20628 14232
rect 20680 14220 20686 14272
rect 20732 14269 20760 14368
rect 22094 14356 22100 14408
rect 22152 14356 22158 14408
rect 22278 14356 22284 14408
rect 22336 14396 22342 14408
rect 23032 14405 23060 14436
rect 22741 14399 22799 14405
rect 22741 14396 22753 14399
rect 22336 14368 22753 14396
rect 22336 14356 22342 14368
rect 22741 14365 22753 14368
rect 22787 14365 22799 14399
rect 22741 14359 22799 14365
rect 23017 14399 23075 14405
rect 23017 14365 23029 14399
rect 23063 14365 23075 14399
rect 23017 14359 23075 14365
rect 21852 14331 21910 14337
rect 21852 14297 21864 14331
rect 21898 14328 21910 14331
rect 22554 14328 22560 14340
rect 21898 14300 22560 14328
rect 21898 14297 21910 14300
rect 21852 14291 21910 14297
rect 22554 14288 22560 14300
rect 22612 14288 22618 14340
rect 23293 14331 23351 14337
rect 23293 14297 23305 14331
rect 23339 14328 23351 14331
rect 23382 14328 23388 14340
rect 23339 14300 23388 14328
rect 23339 14297 23351 14300
rect 23293 14291 23351 14297
rect 23382 14288 23388 14300
rect 23440 14288 23446 14340
rect 20717 14263 20775 14269
rect 20717 14229 20729 14263
rect 20763 14229 20775 14263
rect 20717 14223 20775 14229
rect 21174 14220 21180 14272
rect 21232 14260 21238 14272
rect 22189 14263 22247 14269
rect 22189 14260 22201 14263
rect 21232 14232 22201 14260
rect 21232 14220 21238 14232
rect 22189 14229 22201 14232
rect 22235 14229 22247 14263
rect 22189 14223 22247 14229
rect 1104 14170 23828 14192
rect 1104 14118 2658 14170
rect 2710 14118 2722 14170
rect 2774 14118 2786 14170
rect 2838 14118 2850 14170
rect 2902 14118 2914 14170
rect 2966 14118 2978 14170
rect 3030 14118 8658 14170
rect 8710 14118 8722 14170
rect 8774 14118 8786 14170
rect 8838 14118 8850 14170
rect 8902 14118 8914 14170
rect 8966 14118 8978 14170
rect 9030 14118 14658 14170
rect 14710 14118 14722 14170
rect 14774 14118 14786 14170
rect 14838 14118 14850 14170
rect 14902 14118 14914 14170
rect 14966 14118 14978 14170
rect 15030 14118 20658 14170
rect 20710 14118 20722 14170
rect 20774 14118 20786 14170
rect 20838 14118 20850 14170
rect 20902 14118 20914 14170
rect 20966 14118 20978 14170
rect 21030 14118 23828 14170
rect 1104 14096 23828 14118
rect 1765 14059 1823 14065
rect 1765 14025 1777 14059
rect 1811 14056 1823 14059
rect 6822 14056 6828 14068
rect 1811 14028 6828 14056
rect 1811 14025 1823 14028
rect 1765 14019 1823 14025
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 12986 14056 12992 14068
rect 7852 14028 12992 14056
rect 3694 13988 3700 14000
rect 1596 13960 3700 13988
rect 1596 13929 1624 13960
rect 3694 13948 3700 13960
rect 3752 13948 3758 14000
rect 7592 13991 7650 13997
rect 4080 13960 5672 13988
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13889 1639 13923
rect 1581 13883 1639 13889
rect 1762 13880 1768 13932
rect 1820 13920 1826 13932
rect 2130 13929 2136 13932
rect 1857 13923 1915 13929
rect 1857 13920 1869 13923
rect 1820 13892 1869 13920
rect 1820 13880 1826 13892
rect 1857 13889 1869 13892
rect 1903 13889 1915 13923
rect 2124 13920 2136 13929
rect 2091 13892 2136 13920
rect 1857 13883 1915 13889
rect 2124 13883 2136 13892
rect 2130 13880 2136 13883
rect 2188 13880 2194 13932
rect 3142 13880 3148 13932
rect 3200 13920 3206 13932
rect 3326 13920 3332 13932
rect 3200 13892 3332 13920
rect 3200 13880 3206 13892
rect 3326 13880 3332 13892
rect 3384 13880 3390 13932
rect 3585 13923 3643 13929
rect 3585 13920 3597 13923
rect 3436 13892 3597 13920
rect 3436 13852 3464 13892
rect 3585 13889 3597 13892
rect 3631 13889 3643 13923
rect 3585 13883 3643 13889
rect 3878 13880 3884 13932
rect 3936 13920 3942 13932
rect 4080 13920 4108 13960
rect 5644 13932 5672 13960
rect 7592 13957 7604 13991
rect 7638 13988 7650 13991
rect 7638 13960 7788 13988
rect 7638 13957 7650 13960
rect 7592 13951 7650 13957
rect 3936 13892 4108 13920
rect 3936 13880 3942 13892
rect 4430 13880 4436 13932
rect 4488 13880 4494 13932
rect 5074 13929 5080 13932
rect 5068 13883 5080 13929
rect 5074 13880 5080 13883
rect 5132 13880 5138 13932
rect 5626 13880 5632 13932
rect 5684 13880 5690 13932
rect 3252 13824 3464 13852
rect 4448 13852 4476 13880
rect 4448 13824 4752 13852
rect 3252 13793 3280 13824
rect 4724 13793 4752 13824
rect 4798 13812 4804 13864
rect 4856 13812 4862 13864
rect 7760 13852 7788 13960
rect 7852 13929 7880 14028
rect 12986 14016 12992 14028
rect 13044 14016 13050 14068
rect 13354 14016 13360 14068
rect 13412 14056 13418 14068
rect 13449 14059 13507 14065
rect 13449 14056 13461 14059
rect 13412 14028 13461 14056
rect 13412 14016 13418 14028
rect 13449 14025 13461 14028
rect 13495 14025 13507 14059
rect 13449 14019 13507 14025
rect 14182 14016 14188 14068
rect 14240 14056 14246 14068
rect 15381 14059 15439 14065
rect 15381 14056 15393 14059
rect 14240 14028 15393 14056
rect 14240 14016 14246 14028
rect 15381 14025 15393 14028
rect 15427 14025 15439 14059
rect 15381 14019 15439 14025
rect 16390 14016 16396 14068
rect 16448 14016 16454 14068
rect 16482 14016 16488 14068
rect 16540 14016 16546 14068
rect 16853 14059 16911 14065
rect 16853 14025 16865 14059
rect 16899 14025 16911 14059
rect 16853 14019 16911 14025
rect 16945 14059 17003 14065
rect 16945 14025 16957 14059
rect 16991 14056 17003 14059
rect 17218 14056 17224 14068
rect 16991 14028 17224 14056
rect 16991 14025 17003 14028
rect 16945 14019 17003 14025
rect 9858 13988 9864 14000
rect 7944 13960 8432 13988
rect 7944 13929 7972 13960
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13889 7895 13923
rect 7837 13883 7895 13889
rect 7929 13923 7987 13929
rect 7929 13889 7941 13923
rect 7975 13889 7987 13923
rect 8404 13920 8432 13960
rect 9646 13960 9864 13988
rect 9122 13920 9128 13932
rect 8404 13892 9128 13920
rect 7929 13883 7987 13889
rect 9122 13880 9128 13892
rect 9180 13880 9186 13932
rect 5828 13824 6500 13852
rect 7760 13824 8340 13852
rect 3237 13787 3295 13793
rect 3237 13753 3249 13787
rect 3283 13753 3295 13787
rect 3237 13747 3295 13753
rect 4709 13787 4767 13793
rect 4709 13753 4721 13787
rect 4755 13753 4767 13787
rect 4709 13747 4767 13753
rect 3050 13676 3056 13728
rect 3108 13716 3114 13728
rect 5828 13716 5856 13824
rect 6181 13787 6239 13793
rect 6181 13753 6193 13787
rect 6227 13784 6239 13787
rect 6362 13784 6368 13796
rect 6227 13756 6368 13784
rect 6227 13753 6239 13756
rect 6181 13747 6239 13753
rect 6362 13744 6368 13756
rect 6420 13744 6426 13796
rect 6472 13793 6500 13824
rect 6457 13787 6515 13793
rect 6457 13753 6469 13787
rect 6503 13753 6515 13787
rect 8312 13784 8340 13824
rect 8386 13812 8392 13864
rect 8444 13852 8450 13864
rect 9493 13855 9551 13861
rect 9493 13852 9505 13855
rect 8444 13824 9505 13852
rect 8444 13812 8450 13824
rect 9493 13821 9505 13824
rect 9539 13821 9551 13855
rect 9493 13815 9551 13821
rect 9646 13784 9674 13960
rect 9858 13948 9864 13960
rect 9916 13948 9922 14000
rect 9950 13948 9956 14000
rect 10008 13948 10014 14000
rect 11517 13991 11575 13997
rect 11517 13957 11529 13991
rect 11563 13988 11575 13991
rect 11882 13988 11888 14000
rect 11563 13960 11888 13988
rect 11563 13957 11575 13960
rect 11517 13951 11575 13957
rect 11882 13948 11888 13960
rect 11940 13948 11946 14000
rect 11974 13948 11980 14000
rect 12032 13948 12038 14000
rect 12894 13988 12900 14000
rect 12084 13960 12900 13988
rect 9968 13793 9996 13948
rect 11054 13880 11060 13932
rect 11112 13929 11118 13932
rect 11112 13883 11124 13929
rect 11112 13880 11118 13883
rect 11330 13812 11336 13864
rect 11388 13812 11394 13864
rect 11992 13861 12020 13948
rect 12084 13929 12112 13960
rect 12894 13948 12900 13960
rect 12952 13948 12958 14000
rect 13538 13948 13544 14000
rect 13596 13948 13602 14000
rect 15102 13948 15108 14000
rect 15160 13948 15166 14000
rect 12069 13923 12127 13929
rect 12069 13889 12081 13923
rect 12115 13889 12127 13923
rect 12069 13883 12127 13889
rect 12158 13880 12164 13932
rect 12216 13920 12222 13932
rect 12325 13923 12383 13929
rect 12325 13920 12337 13923
rect 12216 13892 12337 13920
rect 12216 13880 12222 13892
rect 12325 13889 12337 13892
rect 12371 13889 12383 13923
rect 12325 13883 12383 13889
rect 13814 13880 13820 13932
rect 13872 13920 13878 13932
rect 15120 13920 15148 13948
rect 15565 13923 15623 13929
rect 15565 13920 15577 13923
rect 13872 13892 15577 13920
rect 13872 13880 13878 13892
rect 15565 13889 15577 13892
rect 15611 13889 15623 13923
rect 15565 13883 15623 13889
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13920 15991 13923
rect 16408 13920 16436 14016
rect 16868 13988 16896 14019
rect 17218 14016 17224 14028
rect 17276 14016 17282 14068
rect 17678 14016 17684 14068
rect 17736 14016 17742 14068
rect 18138 14016 18144 14068
rect 18196 14016 18202 14068
rect 18230 14016 18236 14068
rect 18288 14016 18294 14068
rect 19334 14016 19340 14068
rect 19392 14056 19398 14068
rect 20625 14059 20683 14065
rect 20625 14056 20637 14059
rect 19392 14028 20637 14056
rect 19392 14016 19398 14028
rect 20625 14025 20637 14028
rect 20671 14025 20683 14059
rect 20625 14019 20683 14025
rect 21266 14016 21272 14068
rect 21324 14016 21330 14068
rect 22094 14016 22100 14068
rect 22152 14056 22158 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 22152 14028 23397 14056
rect 22152 14016 22158 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 23385 14019 23443 14025
rect 18156 13988 18184 14016
rect 16868 13960 18184 13988
rect 15979 13892 16436 13920
rect 16669 13923 16727 13929
rect 15979 13889 15991 13892
rect 15933 13883 15991 13889
rect 16669 13889 16681 13923
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 11977 13855 12035 13861
rect 11977 13821 11989 13855
rect 12023 13821 12035 13855
rect 16684 13852 16712 13883
rect 17034 13880 17040 13932
rect 17092 13920 17098 13932
rect 17497 13923 17555 13929
rect 17497 13920 17509 13923
rect 17092 13892 17509 13920
rect 17092 13880 17098 13892
rect 17497 13889 17509 13892
rect 17543 13889 17555 13923
rect 18248 13920 18276 14016
rect 18506 13948 18512 14000
rect 18564 13988 18570 14000
rect 18794 13991 18852 13997
rect 18794 13988 18806 13991
rect 18564 13960 18806 13988
rect 18564 13948 18570 13960
rect 18794 13957 18806 13960
rect 18840 13957 18852 13991
rect 21284 13988 21312 14016
rect 18794 13951 18852 13957
rect 19076 13960 21312 13988
rect 19076 13929 19104 13960
rect 22646 13948 22652 14000
rect 22704 13948 22710 14000
rect 23198 13948 23204 14000
rect 23256 13948 23262 14000
rect 23290 13948 23296 14000
rect 23348 13948 23354 14000
rect 17497 13883 17555 13889
rect 17604 13892 18276 13920
rect 19061 13923 19119 13929
rect 17604 13852 17632 13892
rect 19061 13889 19073 13923
rect 19107 13889 19119 13923
rect 19978 13920 19984 13932
rect 19061 13883 19119 13889
rect 19168 13892 19984 13920
rect 18046 13852 18052 13864
rect 16684 13824 17632 13852
rect 17972 13824 18052 13852
rect 11977 13815 12035 13821
rect 8312 13756 9674 13784
rect 9953 13787 10011 13793
rect 6457 13747 6515 13753
rect 9953 13753 9965 13787
rect 9999 13753 10011 13787
rect 9953 13747 10011 13753
rect 11606 13744 11612 13796
rect 11664 13784 11670 13796
rect 11793 13787 11851 13793
rect 11793 13784 11805 13787
rect 11664 13756 11805 13784
rect 11664 13744 11670 13756
rect 11793 13753 11805 13756
rect 11839 13753 11851 13787
rect 11793 13747 11851 13753
rect 13814 13744 13820 13796
rect 13872 13784 13878 13796
rect 17126 13784 17132 13796
rect 13872 13756 17132 13784
rect 13872 13744 13878 13756
rect 17126 13744 17132 13756
rect 17184 13784 17190 13796
rect 17972 13784 18000 13824
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 19168 13793 19196 13892
rect 19978 13880 19984 13892
rect 20036 13880 20042 13932
rect 20277 13923 20335 13929
rect 20277 13889 20289 13923
rect 20323 13920 20335 13923
rect 20533 13923 20591 13929
rect 20323 13892 20484 13920
rect 20323 13889 20335 13892
rect 20277 13883 20335 13889
rect 20456 13852 20484 13892
rect 20533 13889 20545 13923
rect 20579 13920 20591 13923
rect 21450 13920 21456 13932
rect 20579 13892 21456 13920
rect 20579 13889 20591 13892
rect 20533 13883 20591 13889
rect 21450 13880 21456 13892
rect 21508 13880 21514 13932
rect 21542 13880 21548 13932
rect 21600 13880 21606 13932
rect 21726 13880 21732 13932
rect 21784 13920 21790 13932
rect 21821 13923 21879 13929
rect 21821 13920 21833 13923
rect 21784 13892 21833 13920
rect 21784 13880 21790 13892
rect 21821 13889 21833 13892
rect 21867 13889 21879 13923
rect 21821 13883 21879 13889
rect 22088 13923 22146 13929
rect 22088 13889 22100 13923
rect 22134 13920 22146 13923
rect 22664 13920 22692 13948
rect 22134 13892 22692 13920
rect 22134 13889 22146 13892
rect 22088 13883 22146 13889
rect 21174 13852 21180 13864
rect 20456 13824 21180 13852
rect 21174 13812 21180 13824
rect 21232 13812 21238 13864
rect 21269 13855 21327 13861
rect 21269 13821 21281 13855
rect 21315 13852 21327 13855
rect 21358 13852 21364 13864
rect 21315 13824 21364 13852
rect 21315 13821 21327 13824
rect 21269 13815 21327 13821
rect 21358 13812 21364 13824
rect 21416 13812 21422 13864
rect 23216 13793 23244 13948
rect 23308 13919 23336 13948
rect 23293 13913 23351 13919
rect 23293 13879 23305 13913
rect 23339 13879 23351 13913
rect 23293 13873 23351 13879
rect 17184 13756 18000 13784
rect 19153 13787 19211 13793
rect 17184 13744 17190 13756
rect 19153 13753 19165 13787
rect 19199 13753 19211 13787
rect 19153 13747 19211 13753
rect 23201 13787 23259 13793
rect 23201 13753 23213 13787
rect 23247 13753 23259 13787
rect 23201 13747 23259 13753
rect 3108 13688 5856 13716
rect 3108 13676 3114 13688
rect 14826 13676 14832 13728
rect 14884 13676 14890 13728
rect 20806 13676 20812 13728
rect 20864 13716 20870 13728
rect 21361 13719 21419 13725
rect 21361 13716 21373 13719
rect 20864 13688 21373 13716
rect 20864 13676 20870 13688
rect 21361 13685 21373 13688
rect 21407 13685 21419 13719
rect 21361 13679 21419 13685
rect 1104 13626 23828 13648
rect 1104 13574 1918 13626
rect 1970 13574 1982 13626
rect 2034 13574 2046 13626
rect 2098 13574 2110 13626
rect 2162 13574 2174 13626
rect 2226 13574 2238 13626
rect 2290 13574 7918 13626
rect 7970 13574 7982 13626
rect 8034 13574 8046 13626
rect 8098 13574 8110 13626
rect 8162 13574 8174 13626
rect 8226 13574 8238 13626
rect 8290 13574 13918 13626
rect 13970 13574 13982 13626
rect 14034 13574 14046 13626
rect 14098 13574 14110 13626
rect 14162 13574 14174 13626
rect 14226 13574 14238 13626
rect 14290 13574 19918 13626
rect 19970 13574 19982 13626
rect 20034 13574 20046 13626
rect 20098 13574 20110 13626
rect 20162 13574 20174 13626
rect 20226 13574 20238 13626
rect 20290 13574 23828 13626
rect 1104 13552 23828 13574
rect 3234 13472 3240 13524
rect 3292 13512 3298 13524
rect 3292 13484 3832 13512
rect 3292 13472 3298 13484
rect 934 13336 940 13388
rect 992 13376 998 13388
rect 1489 13379 1547 13385
rect 1489 13376 1501 13379
rect 992 13348 1501 13376
rect 992 13336 998 13348
rect 1489 13345 1501 13348
rect 1535 13345 1547 13379
rect 1489 13339 1547 13345
rect 2041 13311 2099 13317
rect 2041 13277 2053 13311
rect 2087 13308 2099 13311
rect 3050 13308 3056 13320
rect 2087 13280 3056 13308
rect 2087 13277 2099 13280
rect 2041 13271 2099 13277
rect 3050 13268 3056 13280
rect 3108 13268 3114 13320
rect 3510 13268 3516 13320
rect 3568 13308 3574 13320
rect 3804 13317 3832 13484
rect 3896 13484 9168 13512
rect 3896 13453 3924 13484
rect 3881 13447 3939 13453
rect 3881 13413 3893 13447
rect 3927 13413 3939 13447
rect 3881 13407 3939 13413
rect 7006 13404 7012 13456
rect 7064 13444 7070 13456
rect 7285 13447 7343 13453
rect 7285 13444 7297 13447
rect 7064 13416 7297 13444
rect 7064 13404 7070 13416
rect 7285 13413 7297 13416
rect 7331 13413 7343 13447
rect 9140 13444 9168 13484
rect 10778 13472 10784 13524
rect 10836 13472 10842 13524
rect 12894 13472 12900 13524
rect 12952 13472 12958 13524
rect 12986 13472 12992 13524
rect 13044 13512 13050 13524
rect 13541 13515 13599 13521
rect 13541 13512 13553 13515
rect 13044 13484 13553 13512
rect 13044 13472 13050 13484
rect 13541 13481 13553 13484
rect 13587 13481 13599 13515
rect 14366 13512 14372 13524
rect 13541 13475 13599 13481
rect 13924 13484 14372 13512
rect 9674 13444 9680 13456
rect 9140 13416 9680 13444
rect 7285 13407 7343 13413
rect 9674 13404 9680 13416
rect 9732 13404 9738 13456
rect 12912 13444 12940 13472
rect 13817 13447 13875 13453
rect 13817 13444 13829 13447
rect 12912 13416 13829 13444
rect 13817 13413 13829 13416
rect 13863 13413 13875 13447
rect 13817 13407 13875 13413
rect 4062 13336 4068 13388
rect 4120 13336 4126 13388
rect 13170 13336 13176 13388
rect 13228 13336 13234 13388
rect 3605 13311 3663 13317
rect 3605 13308 3617 13311
rect 3568 13280 3617 13308
rect 3568 13268 3574 13280
rect 3605 13277 3617 13280
rect 3651 13277 3663 13311
rect 3605 13271 3663 13277
rect 3789 13311 3847 13317
rect 3789 13277 3801 13311
rect 3835 13308 3847 13311
rect 5537 13311 5595 13317
rect 3835 13280 4476 13308
rect 3835 13277 3847 13280
rect 3789 13271 3847 13277
rect 3234 13240 3240 13252
rect 2746 13212 3240 13240
rect 2225 13175 2283 13181
rect 2225 13141 2237 13175
rect 2271 13172 2283 13175
rect 2746 13172 2774 13212
rect 3234 13200 3240 13212
rect 3292 13200 3298 13252
rect 3326 13200 3332 13252
rect 3384 13249 3390 13252
rect 4338 13249 4344 13252
rect 3384 13203 3396 13249
rect 4332 13203 4344 13249
rect 3384 13200 3390 13203
rect 4338 13200 4344 13203
rect 4396 13200 4402 13252
rect 4448 13240 4476 13280
rect 5537 13277 5549 13311
rect 5583 13308 5595 13311
rect 6638 13308 6644 13320
rect 5583 13280 6644 13308
rect 5583 13277 5595 13280
rect 5537 13271 5595 13277
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 10689 13311 10747 13317
rect 10689 13277 10701 13311
rect 10735 13308 10747 13311
rect 11146 13308 11152 13320
rect 10735 13280 11152 13308
rect 10735 13277 10747 13280
rect 10689 13271 10747 13277
rect 11146 13268 11152 13280
rect 11204 13268 11210 13320
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 11333 13311 11391 13317
rect 11333 13308 11345 13311
rect 11296 13280 11345 13308
rect 11296 13268 11302 13280
rect 11333 13277 11345 13280
rect 11379 13277 11391 13311
rect 11333 13271 11391 13277
rect 11606 13268 11612 13320
rect 11664 13268 11670 13320
rect 11882 13268 11888 13320
rect 11940 13268 11946 13320
rect 13446 13268 13452 13320
rect 13504 13268 13510 13320
rect 13924 13317 13952 13484
rect 14366 13472 14372 13484
rect 14424 13512 14430 13524
rect 14424 13484 15884 13512
rect 14424 13472 14430 13484
rect 14277 13447 14335 13453
rect 14277 13413 14289 13447
rect 14323 13444 14335 13447
rect 15378 13444 15384 13456
rect 14323 13416 15384 13444
rect 14323 13413 14335 13416
rect 14277 13407 14335 13413
rect 15378 13404 15384 13416
rect 15436 13404 15442 13456
rect 15856 13444 15884 13484
rect 15930 13472 15936 13524
rect 15988 13512 15994 13524
rect 16761 13515 16819 13521
rect 16761 13512 16773 13515
rect 15988 13484 16773 13512
rect 15988 13472 15994 13484
rect 16761 13481 16773 13484
rect 16807 13481 16819 13515
rect 16761 13475 16819 13481
rect 18693 13515 18751 13521
rect 18693 13481 18705 13515
rect 18739 13512 18751 13515
rect 19886 13512 19892 13524
rect 18739 13484 19892 13512
rect 18739 13481 18751 13484
rect 18693 13475 18751 13481
rect 19886 13472 19892 13484
rect 19944 13472 19950 13524
rect 22097 13515 22155 13521
rect 22097 13481 22109 13515
rect 22143 13512 22155 13515
rect 22186 13512 22192 13524
rect 22143 13484 22192 13512
rect 22143 13481 22155 13484
rect 22097 13475 22155 13481
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 16390 13444 16396 13456
rect 15856 13416 16396 13444
rect 16390 13404 16396 13416
rect 16448 13404 16454 13456
rect 14826 13376 14832 13388
rect 14384 13348 14832 13376
rect 14384 13317 14412 13348
rect 14826 13336 14832 13348
rect 14884 13336 14890 13388
rect 23382 13336 23388 13388
rect 23440 13336 23446 13388
rect 13909 13311 13967 13317
rect 13909 13277 13921 13311
rect 13955 13277 13967 13311
rect 13909 13271 13967 13277
rect 14093 13311 14151 13317
rect 14093 13277 14105 13311
rect 14139 13308 14151 13311
rect 14369 13311 14427 13317
rect 14369 13308 14381 13311
rect 14139 13280 14381 13308
rect 14139 13277 14151 13280
rect 14093 13271 14151 13277
rect 14369 13277 14381 13280
rect 14415 13277 14427 13311
rect 14369 13271 14427 13277
rect 14737 13311 14795 13317
rect 14737 13277 14749 13311
rect 14783 13308 14795 13311
rect 17034 13308 17040 13320
rect 14783 13280 17040 13308
rect 14783 13277 14795 13280
rect 14737 13271 14795 13277
rect 5810 13249 5816 13252
rect 4448 13212 5580 13240
rect 2271 13144 2774 13172
rect 2271 13141 2283 13144
rect 2225 13135 2283 13141
rect 3142 13132 3148 13184
rect 3200 13172 3206 13184
rect 5350 13172 5356 13184
rect 3200 13144 5356 13172
rect 3200 13132 3206 13144
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 5442 13132 5448 13184
rect 5500 13132 5506 13184
rect 5552 13172 5580 13212
rect 5804 13203 5816 13249
rect 5810 13200 5816 13203
rect 5868 13200 5874 13252
rect 8386 13240 8392 13252
rect 6380 13212 8392 13240
rect 6380 13172 6408 13212
rect 8386 13200 8392 13212
rect 8444 13200 8450 13252
rect 8757 13243 8815 13249
rect 8757 13209 8769 13243
rect 8803 13209 8815 13243
rect 8757 13203 8815 13209
rect 5552 13144 6408 13172
rect 6917 13175 6975 13181
rect 6917 13141 6929 13175
rect 6963 13172 6975 13175
rect 7190 13172 7196 13184
rect 6963 13144 7196 13172
rect 6963 13141 6975 13144
rect 6917 13135 6975 13141
rect 7190 13132 7196 13144
rect 7248 13132 7254 13184
rect 8772 13172 8800 13203
rect 9030 13200 9036 13252
rect 9088 13240 9094 13252
rect 9088 13212 9444 13240
rect 9088 13200 9094 13212
rect 9306 13172 9312 13184
rect 8772 13144 9312 13172
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 9416 13181 9444 13212
rect 9401 13175 9459 13181
rect 9401 13141 9413 13175
rect 9447 13172 9459 13175
rect 9490 13172 9496 13184
rect 9447 13144 9496 13172
rect 9447 13141 9459 13144
rect 9401 13135 9459 13141
rect 9490 13132 9496 13144
rect 9548 13132 9554 13184
rect 11146 13132 11152 13184
rect 11204 13172 11210 13184
rect 11900 13172 11928 13268
rect 13814 13200 13820 13252
rect 13872 13240 13878 13252
rect 14108 13240 14136 13271
rect 17034 13268 17040 13280
rect 17092 13268 17098 13320
rect 17310 13268 17316 13320
rect 17368 13268 17374 13320
rect 18046 13308 18052 13320
rect 17512 13280 18052 13308
rect 13872 13212 14136 13240
rect 13872 13200 13878 13212
rect 15470 13200 15476 13252
rect 15528 13200 15534 13252
rect 11204 13144 11928 13172
rect 14553 13175 14611 13181
rect 11204 13132 11210 13144
rect 14553 13141 14565 13175
rect 14599 13172 14611 13175
rect 15286 13172 15292 13184
rect 14599 13144 15292 13172
rect 14599 13141 14611 13144
rect 14553 13135 14611 13141
rect 15286 13132 15292 13144
rect 15344 13132 15350 13184
rect 15381 13175 15439 13181
rect 15381 13141 15393 13175
rect 15427 13172 15439 13175
rect 17512 13172 17540 13280
rect 18046 13268 18052 13280
rect 18104 13268 18110 13320
rect 18969 13311 19027 13317
rect 18969 13277 18981 13311
rect 19015 13277 19027 13311
rect 18969 13271 19027 13277
rect 17580 13243 17638 13249
rect 17580 13209 17592 13243
rect 17626 13240 17638 13243
rect 17626 13212 17908 13240
rect 17626 13209 17638 13212
rect 17580 13203 17638 13209
rect 15427 13144 17540 13172
rect 17880 13172 17908 13212
rect 17954 13200 17960 13252
rect 18012 13240 18018 13252
rect 18984 13240 19012 13271
rect 19334 13268 19340 13320
rect 19392 13308 19398 13320
rect 20625 13311 20683 13317
rect 20625 13308 20637 13311
rect 19392 13280 20637 13308
rect 19392 13268 19398 13280
rect 20625 13277 20637 13280
rect 20671 13277 20683 13311
rect 20625 13271 20683 13277
rect 20717 13311 20775 13317
rect 20717 13277 20729 13311
rect 20763 13308 20775 13311
rect 21542 13308 21548 13320
rect 20763 13280 21548 13308
rect 20763 13277 20775 13280
rect 20717 13271 20775 13277
rect 21542 13268 21548 13280
rect 21600 13268 21606 13320
rect 21818 13268 21824 13320
rect 21876 13308 21882 13320
rect 22189 13311 22247 13317
rect 22189 13308 22201 13311
rect 21876 13280 22201 13308
rect 21876 13268 21882 13280
rect 22189 13277 22201 13280
rect 22235 13277 22247 13311
rect 22189 13271 22247 13277
rect 22370 13268 22376 13320
rect 22428 13308 22434 13320
rect 22833 13311 22891 13317
rect 22833 13308 22845 13311
rect 22428 13280 22845 13308
rect 22428 13268 22434 13280
rect 22833 13277 22845 13280
rect 22879 13277 22891 13311
rect 22833 13271 22891 13277
rect 18012 13212 19012 13240
rect 20380 13243 20438 13249
rect 18012 13200 18018 13212
rect 20380 13209 20392 13243
rect 20426 13240 20438 13243
rect 20806 13240 20812 13252
rect 20426 13212 20812 13240
rect 20426 13209 20438 13212
rect 20380 13203 20438 13209
rect 20806 13200 20812 13212
rect 20864 13200 20870 13252
rect 20984 13243 21042 13249
rect 20984 13209 20996 13243
rect 21030 13209 21042 13243
rect 20984 13203 21042 13209
rect 22465 13243 22523 13249
rect 22465 13209 22477 13243
rect 22511 13240 22523 13243
rect 23382 13240 23388 13252
rect 22511 13212 23388 13240
rect 22511 13209 22523 13212
rect 22465 13203 22523 13209
rect 18138 13172 18144 13184
rect 17880 13144 18144 13172
rect 15427 13141 15439 13144
rect 15381 13135 15439 13141
rect 18138 13132 18144 13144
rect 18196 13132 18202 13184
rect 18874 13132 18880 13184
rect 18932 13132 18938 13184
rect 19242 13132 19248 13184
rect 19300 13132 19306 13184
rect 19978 13132 19984 13184
rect 20036 13172 20042 13184
rect 21008 13172 21036 13203
rect 23382 13200 23388 13212
rect 23440 13200 23446 13252
rect 20036 13144 21036 13172
rect 20036 13132 20042 13144
rect 1104 13082 23828 13104
rect 1104 13030 2658 13082
rect 2710 13030 2722 13082
rect 2774 13030 2786 13082
rect 2838 13030 2850 13082
rect 2902 13030 2914 13082
rect 2966 13030 2978 13082
rect 3030 13030 8658 13082
rect 8710 13030 8722 13082
rect 8774 13030 8786 13082
rect 8838 13030 8850 13082
rect 8902 13030 8914 13082
rect 8966 13030 8978 13082
rect 9030 13030 14658 13082
rect 14710 13030 14722 13082
rect 14774 13030 14786 13082
rect 14838 13030 14850 13082
rect 14902 13030 14914 13082
rect 14966 13030 14978 13082
rect 15030 13030 20658 13082
rect 20710 13030 20722 13082
rect 20774 13030 20786 13082
rect 20838 13030 20850 13082
rect 20902 13030 20914 13082
rect 20966 13030 20978 13082
rect 21030 13030 23828 13082
rect 1104 13008 23828 13030
rect 1673 12971 1731 12977
rect 1673 12937 1685 12971
rect 1719 12968 1731 12971
rect 4798 12968 4804 12980
rect 1719 12940 4804 12968
rect 1719 12937 1731 12940
rect 1673 12931 1731 12937
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 5350 12928 5356 12980
rect 5408 12968 5414 12980
rect 6457 12971 6515 12977
rect 5408 12940 6408 12968
rect 5408 12928 5414 12940
rect 3142 12900 3148 12912
rect 2746 12872 3148 12900
rect 1765 12835 1823 12841
rect 1765 12801 1777 12835
rect 1811 12832 1823 12835
rect 2746 12832 2774 12872
rect 3142 12860 3148 12872
rect 3200 12860 3206 12912
rect 4706 12900 4712 12912
rect 3344 12872 4712 12900
rect 1811 12804 2774 12832
rect 1811 12801 1823 12804
rect 1765 12795 1823 12801
rect 2958 12792 2964 12844
rect 3016 12841 3022 12844
rect 3344 12841 3372 12872
rect 4706 12860 4712 12872
rect 4764 12860 4770 12912
rect 3016 12835 3039 12841
rect 3027 12801 3039 12835
rect 3016 12795 3039 12801
rect 3237 12835 3295 12841
rect 3237 12801 3249 12835
rect 3283 12832 3295 12835
rect 3329 12835 3387 12841
rect 3329 12832 3341 12835
rect 3283 12804 3341 12832
rect 3283 12801 3295 12804
rect 3237 12795 3295 12801
rect 3329 12801 3341 12804
rect 3375 12801 3387 12835
rect 3329 12795 3387 12801
rect 3016 12792 3022 12795
rect 3418 12792 3424 12844
rect 3476 12832 3482 12844
rect 3585 12835 3643 12841
rect 3585 12832 3597 12835
rect 3476 12804 3597 12832
rect 3476 12792 3482 12804
rect 3585 12801 3597 12804
rect 3631 12801 3643 12835
rect 3585 12795 3643 12801
rect 4890 12792 4896 12844
rect 4948 12832 4954 12844
rect 6380 12841 6408 12940
rect 6457 12937 6469 12971
rect 6503 12968 6515 12971
rect 11330 12968 11336 12980
rect 6503 12940 11336 12968
rect 6503 12937 6515 12940
rect 6457 12931 6515 12937
rect 11330 12928 11336 12940
rect 11388 12928 11394 12980
rect 12802 12968 12808 12980
rect 12406 12940 12808 12968
rect 6733 12903 6791 12909
rect 6733 12869 6745 12903
rect 6779 12900 6791 12903
rect 10873 12903 10931 12909
rect 6779 12872 10824 12900
rect 6779 12869 6791 12872
rect 6733 12863 6791 12869
rect 5057 12835 5115 12841
rect 5057 12832 5069 12835
rect 4948 12804 5069 12832
rect 4948 12792 4954 12804
rect 5057 12801 5069 12804
rect 5103 12801 5115 12835
rect 5057 12795 5115 12801
rect 6365 12835 6423 12841
rect 6365 12801 6377 12835
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 4801 12767 4859 12773
rect 4801 12764 4813 12767
rect 4540 12736 4813 12764
rect 1762 12588 1768 12640
rect 1820 12628 1826 12640
rect 1857 12631 1915 12637
rect 1857 12628 1869 12631
rect 1820 12600 1869 12628
rect 1820 12588 1826 12600
rect 1857 12597 1869 12600
rect 1903 12597 1915 12631
rect 1857 12591 1915 12597
rect 3510 12588 3516 12640
rect 3568 12628 3574 12640
rect 4540 12628 4568 12736
rect 4801 12733 4813 12736
rect 4847 12733 4859 12767
rect 6380 12764 6408 12795
rect 6822 12792 6828 12844
rect 6880 12792 6886 12844
rect 7009 12835 7067 12841
rect 7009 12801 7021 12835
rect 7055 12832 7067 12835
rect 7190 12832 7196 12844
rect 7055 12804 7196 12832
rect 7055 12801 7067 12804
rect 7009 12795 7067 12801
rect 7190 12792 7196 12804
rect 7248 12792 7254 12844
rect 7650 12792 7656 12844
rect 7708 12792 7714 12844
rect 7909 12835 7967 12841
rect 7909 12832 7921 12835
rect 7760 12804 7921 12832
rect 6730 12764 6736 12776
rect 6380 12736 6736 12764
rect 4801 12727 4859 12733
rect 6730 12724 6736 12736
rect 6788 12724 6794 12776
rect 7760 12764 7788 12804
rect 7909 12801 7921 12804
rect 7955 12801 7967 12835
rect 7909 12795 7967 12801
rect 8386 12792 8392 12844
rect 8444 12832 8450 12844
rect 8444 12804 9904 12832
rect 8444 12792 8450 12804
rect 7484 12736 7788 12764
rect 4614 12656 4620 12708
rect 4672 12656 4678 12708
rect 3568 12600 4568 12628
rect 4632 12628 4660 12656
rect 7484 12640 7512 12736
rect 7650 12656 7656 12708
rect 7708 12656 7714 12708
rect 9766 12696 9772 12708
rect 8680 12668 9772 12696
rect 4709 12631 4767 12637
rect 4709 12628 4721 12631
rect 4632 12600 4721 12628
rect 3568 12588 3574 12600
rect 4709 12597 4721 12600
rect 4755 12597 4767 12631
rect 4709 12591 4767 12597
rect 6178 12588 6184 12640
rect 6236 12588 6242 12640
rect 7466 12588 7472 12640
rect 7524 12588 7530 12640
rect 7558 12588 7564 12640
rect 7616 12588 7622 12640
rect 7668 12628 7696 12656
rect 8680 12628 8708 12668
rect 9766 12656 9772 12668
rect 9824 12656 9830 12708
rect 9876 12696 9904 12804
rect 10796 12764 10824 12872
rect 10873 12869 10885 12903
rect 10919 12900 10931 12903
rect 12406 12900 12434 12940
rect 12802 12928 12808 12940
rect 12860 12928 12866 12980
rect 13817 12971 13875 12977
rect 13817 12937 13829 12971
rect 13863 12968 13875 12971
rect 16850 12968 16856 12980
rect 13863 12940 16856 12968
rect 13863 12937 13875 12940
rect 13817 12931 13875 12937
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 17034 12928 17040 12980
rect 17092 12968 17098 12980
rect 18325 12971 18383 12977
rect 18325 12968 18337 12971
rect 17092 12940 18337 12968
rect 17092 12928 17098 12940
rect 18325 12937 18337 12940
rect 18371 12937 18383 12971
rect 18325 12931 18383 12937
rect 18874 12928 18880 12980
rect 18932 12928 18938 12980
rect 19242 12928 19248 12980
rect 19300 12928 19306 12980
rect 19794 12928 19800 12980
rect 19852 12928 19858 12980
rect 15194 12900 15200 12912
rect 10919 12872 12434 12900
rect 13556 12872 15200 12900
rect 10919 12869 10931 12872
rect 10873 12863 10931 12869
rect 11330 12792 11336 12844
rect 11388 12792 11394 12844
rect 11514 12792 11520 12844
rect 11572 12792 11578 12844
rect 13556 12841 13584 12872
rect 15194 12860 15200 12872
rect 15252 12860 15258 12912
rect 18892 12900 18920 12928
rect 15856 12872 18920 12900
rect 13541 12835 13599 12841
rect 13541 12801 13553 12835
rect 13587 12801 13599 12835
rect 13541 12795 13599 12801
rect 13630 12792 13636 12844
rect 13688 12792 13694 12844
rect 13906 12792 13912 12844
rect 13964 12792 13970 12844
rect 15102 12832 15108 12844
rect 14752 12804 15108 12832
rect 11606 12764 11612 12776
rect 10796 12736 11612 12764
rect 11606 12724 11612 12736
rect 11664 12724 11670 12776
rect 11422 12696 11428 12708
rect 9876 12668 11428 12696
rect 7668 12600 8708 12628
rect 9033 12631 9091 12637
rect 9033 12597 9045 12631
rect 9079 12628 9091 12631
rect 9398 12628 9404 12640
rect 9079 12600 9404 12628
rect 9079 12597 9091 12600
rect 9033 12591 9091 12597
rect 9398 12588 9404 12600
rect 9456 12588 9462 12640
rect 9585 12631 9643 12637
rect 9585 12597 9597 12631
rect 9631 12628 9643 12631
rect 9876 12628 9904 12668
rect 11422 12656 11428 12668
rect 11480 12656 11486 12708
rect 14274 12656 14280 12708
rect 14332 12656 14338 12708
rect 14461 12699 14519 12705
rect 14461 12665 14473 12699
rect 14507 12696 14519 12699
rect 14752 12696 14780 12804
rect 15102 12792 15108 12804
rect 15160 12792 15166 12844
rect 15856 12841 15884 12872
rect 15585 12835 15643 12841
rect 15585 12801 15597 12835
rect 15631 12832 15643 12835
rect 15841 12835 15899 12841
rect 15631 12804 15792 12832
rect 15631 12801 15643 12804
rect 15585 12795 15643 12801
rect 15764 12764 15792 12804
rect 15841 12801 15853 12835
rect 15887 12801 15899 12835
rect 15841 12795 15899 12801
rect 15933 12835 15991 12841
rect 15933 12801 15945 12835
rect 15979 12832 15991 12835
rect 16853 12835 16911 12841
rect 15979 12804 16804 12832
rect 15979 12801 15991 12804
rect 15933 12795 15991 12801
rect 16666 12764 16672 12776
rect 15764 12736 15884 12764
rect 14507 12668 14780 12696
rect 15856 12696 15884 12736
rect 16132 12736 16672 12764
rect 16132 12696 16160 12736
rect 16666 12724 16672 12736
rect 16724 12724 16730 12776
rect 15856 12668 16160 12696
rect 14507 12665 14519 12668
rect 14461 12659 14519 12665
rect 16206 12656 16212 12708
rect 16264 12656 16270 12708
rect 16776 12696 16804 12804
rect 16853 12801 16865 12835
rect 16899 12832 16911 12835
rect 16942 12832 16948 12844
rect 16899 12804 16948 12832
rect 16899 12801 16911 12804
rect 16853 12795 16911 12801
rect 16942 12792 16948 12804
rect 17000 12792 17006 12844
rect 17120 12835 17178 12841
rect 17120 12801 17132 12835
rect 17166 12832 17178 12835
rect 19260 12832 19288 12928
rect 21634 12900 21640 12912
rect 19720 12872 21640 12900
rect 17166 12804 19288 12832
rect 19449 12835 19507 12841
rect 17166 12801 17178 12804
rect 17120 12795 17178 12801
rect 19449 12801 19461 12835
rect 19495 12832 19507 12835
rect 19610 12832 19616 12844
rect 19495 12804 19616 12832
rect 19495 12801 19507 12804
rect 19449 12795 19507 12801
rect 19610 12792 19616 12804
rect 19668 12792 19674 12844
rect 19720 12773 19748 12872
rect 21634 12860 21640 12872
rect 21692 12860 21698 12912
rect 22088 12903 22146 12909
rect 22088 12869 22100 12903
rect 22134 12900 22146 12903
rect 22186 12900 22192 12912
rect 22134 12872 22192 12900
rect 22134 12869 22146 12872
rect 22088 12863 22146 12869
rect 22186 12860 22192 12872
rect 22244 12860 22250 12912
rect 19886 12792 19892 12844
rect 19944 12832 19950 12844
rect 20910 12835 20968 12841
rect 20910 12832 20922 12835
rect 19944 12804 20922 12832
rect 19944 12792 19950 12804
rect 20910 12801 20922 12804
rect 20956 12801 20968 12835
rect 20910 12795 20968 12801
rect 21082 12792 21088 12844
rect 21140 12832 21146 12844
rect 21358 12832 21364 12844
rect 21140 12804 21364 12832
rect 21140 12792 21146 12804
rect 21358 12792 21364 12804
rect 21416 12832 21422 12844
rect 21453 12835 21511 12841
rect 21453 12832 21465 12835
rect 21416 12804 21465 12832
rect 21416 12792 21422 12804
rect 21453 12801 21465 12804
rect 21499 12801 21511 12835
rect 21453 12795 21511 12801
rect 22370 12792 22376 12844
rect 22428 12832 22434 12844
rect 23293 12835 23351 12841
rect 23293 12832 23305 12835
rect 22428 12804 23305 12832
rect 22428 12792 22434 12804
rect 23293 12801 23305 12804
rect 23339 12801 23351 12835
rect 23293 12795 23351 12801
rect 19705 12767 19763 12773
rect 19705 12733 19717 12767
rect 19751 12733 19763 12767
rect 19705 12727 19763 12733
rect 19978 12724 19984 12776
rect 20036 12724 20042 12776
rect 21177 12767 21235 12773
rect 21177 12733 21189 12767
rect 21223 12764 21235 12767
rect 21726 12764 21732 12776
rect 21223 12736 21732 12764
rect 21223 12733 21235 12736
rect 21177 12727 21235 12733
rect 21726 12724 21732 12736
rect 21784 12724 21790 12776
rect 21821 12767 21879 12773
rect 21821 12733 21833 12767
rect 21867 12733 21879 12767
rect 21821 12727 21879 12733
rect 16850 12696 16856 12708
rect 16776 12668 16856 12696
rect 16850 12656 16856 12668
rect 16908 12656 16914 12708
rect 18233 12699 18291 12705
rect 18233 12665 18245 12699
rect 18279 12696 18291 12699
rect 18279 12668 18828 12696
rect 18279 12665 18291 12668
rect 18233 12659 18291 12665
rect 9631 12600 9904 12628
rect 9631 12597 9643 12600
rect 9585 12591 9643 12597
rect 11146 12588 11152 12640
rect 11204 12588 11210 12640
rect 11330 12588 11336 12640
rect 11388 12628 11394 12640
rect 11790 12628 11796 12640
rect 11388 12600 11796 12628
rect 11388 12588 11394 12600
rect 11790 12588 11796 12600
rect 11848 12588 11854 12640
rect 13449 12631 13507 12637
rect 13449 12597 13461 12631
rect 13495 12628 13507 12631
rect 13722 12628 13728 12640
rect 13495 12600 13728 12628
rect 13495 12597 13507 12600
rect 13449 12591 13507 12597
rect 13722 12588 13728 12600
rect 13780 12588 13786 12640
rect 14366 12588 14372 12640
rect 14424 12588 14430 12640
rect 16393 12631 16451 12637
rect 16393 12597 16405 12631
rect 16439 12628 16451 12631
rect 17586 12628 17592 12640
rect 16439 12600 17592 12628
rect 16439 12597 16451 12600
rect 16393 12591 16451 12597
rect 17586 12588 17592 12600
rect 17644 12588 17650 12640
rect 18800 12628 18828 12668
rect 19996 12628 20024 12724
rect 18800 12600 20024 12628
rect 20438 12588 20444 12640
rect 20496 12628 20502 12640
rect 21361 12631 21419 12637
rect 21361 12628 21373 12631
rect 20496 12600 21373 12628
rect 20496 12588 20502 12600
rect 21361 12597 21373 12600
rect 21407 12597 21419 12631
rect 21361 12591 21419 12597
rect 21726 12588 21732 12640
rect 21784 12628 21790 12640
rect 21836 12628 21864 12727
rect 22830 12724 22836 12776
rect 22888 12764 22894 12776
rect 23385 12767 23443 12773
rect 23385 12764 23397 12767
rect 22888 12736 23397 12764
rect 22888 12724 22894 12736
rect 23385 12733 23397 12736
rect 23431 12733 23443 12767
rect 23385 12727 23443 12733
rect 21784 12600 21864 12628
rect 21784 12588 21790 12600
rect 22554 12588 22560 12640
rect 22612 12628 22618 12640
rect 23201 12631 23259 12637
rect 23201 12628 23213 12631
rect 22612 12600 23213 12628
rect 22612 12588 22618 12600
rect 23201 12597 23213 12600
rect 23247 12597 23259 12631
rect 23201 12591 23259 12597
rect 1104 12538 23828 12560
rect 1104 12486 1918 12538
rect 1970 12486 1982 12538
rect 2034 12486 2046 12538
rect 2098 12486 2110 12538
rect 2162 12486 2174 12538
rect 2226 12486 2238 12538
rect 2290 12486 7918 12538
rect 7970 12486 7982 12538
rect 8034 12486 8046 12538
rect 8098 12486 8110 12538
rect 8162 12486 8174 12538
rect 8226 12486 8238 12538
rect 8290 12486 13918 12538
rect 13970 12486 13982 12538
rect 14034 12486 14046 12538
rect 14098 12486 14110 12538
rect 14162 12486 14174 12538
rect 14226 12486 14238 12538
rect 14290 12486 19918 12538
rect 19970 12486 19982 12538
rect 20034 12486 20046 12538
rect 20098 12486 20110 12538
rect 20162 12486 20174 12538
rect 20226 12486 20238 12538
rect 20290 12486 23828 12538
rect 1104 12464 23828 12486
rect 3326 12384 3332 12436
rect 3384 12424 3390 12436
rect 3605 12427 3663 12433
rect 3605 12424 3617 12427
rect 3384 12396 3617 12424
rect 3384 12384 3390 12396
rect 3605 12393 3617 12396
rect 3651 12393 3663 12427
rect 3605 12387 3663 12393
rect 7650 12384 7656 12436
rect 7708 12424 7714 12436
rect 7708 12396 9720 12424
rect 7708 12384 7714 12396
rect 9692 12356 9720 12396
rect 10226 12384 10232 12436
rect 10284 12424 10290 12436
rect 13446 12424 13452 12436
rect 10284 12396 13452 12424
rect 10284 12384 10290 12396
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 13538 12384 13544 12436
rect 13596 12384 13602 12436
rect 13725 12427 13783 12433
rect 13725 12393 13737 12427
rect 13771 12424 13783 12427
rect 14550 12424 14556 12436
rect 13771 12396 14556 12424
rect 13771 12393 13783 12396
rect 13725 12387 13783 12393
rect 14550 12384 14556 12396
rect 14608 12384 14614 12436
rect 15286 12384 15292 12436
rect 15344 12424 15350 12436
rect 22649 12427 22707 12433
rect 15344 12396 19288 12424
rect 15344 12384 15350 12396
rect 11609 12359 11667 12365
rect 11609 12356 11621 12359
rect 9692 12328 11621 12356
rect 11609 12325 11621 12328
rect 11655 12325 11667 12359
rect 11609 12319 11667 12325
rect 12069 12359 12127 12365
rect 12069 12325 12081 12359
rect 12115 12356 12127 12359
rect 12342 12356 12348 12368
rect 12115 12328 12348 12356
rect 12115 12325 12127 12328
rect 12069 12319 12127 12325
rect 12342 12316 12348 12328
rect 12400 12316 12406 12368
rect 1394 12248 1400 12300
rect 1452 12288 1458 12300
rect 2225 12291 2283 12297
rect 2225 12288 2237 12291
rect 1452 12260 2237 12288
rect 1452 12248 1458 12260
rect 2225 12257 2237 12260
rect 2271 12257 2283 12291
rect 2225 12251 2283 12257
rect 4338 12248 4344 12300
rect 4396 12248 4402 12300
rect 8757 12291 8815 12297
rect 8757 12257 8769 12291
rect 8803 12288 8815 12291
rect 9398 12288 9404 12300
rect 8803 12260 9404 12288
rect 8803 12257 8815 12260
rect 8757 12251 8815 12257
rect 9398 12248 9404 12260
rect 9456 12248 9462 12300
rect 13446 12248 13452 12300
rect 13504 12248 13510 12300
rect 934 12180 940 12232
rect 992 12220 998 12232
rect 1489 12223 1547 12229
rect 1489 12220 1501 12223
rect 992 12192 1501 12220
rect 992 12180 998 12192
rect 1489 12189 1501 12192
rect 1535 12189 1547 12223
rect 1489 12183 1547 12189
rect 2041 12223 2099 12229
rect 2041 12189 2053 12223
rect 2087 12189 2099 12223
rect 2041 12183 2099 12189
rect 2056 12084 2084 12183
rect 3326 12180 3332 12232
rect 3384 12220 3390 12232
rect 7285 12223 7343 12229
rect 3384 12192 4936 12220
rect 3384 12180 3390 12192
rect 4908 12164 4936 12192
rect 7285 12189 7297 12223
rect 7331 12189 7343 12223
rect 7285 12183 7343 12189
rect 8501 12223 8559 12229
rect 8501 12189 8513 12223
rect 8547 12220 8559 12223
rect 8547 12192 8892 12220
rect 8547 12189 8559 12192
rect 8501 12183 8559 12189
rect 2492 12155 2550 12161
rect 2492 12121 2504 12155
rect 2538 12152 2550 12155
rect 3970 12152 3976 12164
rect 2538 12124 3976 12152
rect 2538 12121 2550 12124
rect 2492 12115 2550 12121
rect 3970 12112 3976 12124
rect 4028 12112 4034 12164
rect 4154 12112 4160 12164
rect 4212 12152 4218 12164
rect 4586 12155 4644 12161
rect 4586 12152 4598 12155
rect 4212 12124 4598 12152
rect 4212 12112 4218 12124
rect 4586 12121 4598 12124
rect 4632 12121 4644 12155
rect 4586 12115 4644 12121
rect 4890 12112 4896 12164
rect 4948 12112 4954 12164
rect 7040 12155 7098 12161
rect 7040 12121 7052 12155
rect 7086 12152 7098 12155
rect 7190 12152 7196 12164
rect 7086 12124 7196 12152
rect 7086 12121 7098 12124
rect 7040 12115 7098 12121
rect 7190 12112 7196 12124
rect 7248 12112 7254 12164
rect 7300 12152 7328 12183
rect 8386 12152 8392 12164
rect 7300 12124 8392 12152
rect 8386 12112 8392 12124
rect 8444 12112 8450 12164
rect 8864 12152 8892 12192
rect 8938 12180 8944 12232
rect 8996 12180 9002 12232
rect 9858 12180 9864 12232
rect 9916 12220 9922 12232
rect 10781 12223 10839 12229
rect 10781 12220 10793 12223
rect 9916 12192 10793 12220
rect 9916 12180 9922 12192
rect 10781 12189 10793 12192
rect 10827 12189 10839 12223
rect 10781 12183 10839 12189
rect 11333 12223 11391 12229
rect 11333 12189 11345 12223
rect 11379 12189 11391 12223
rect 11333 12183 11391 12189
rect 13193 12223 13251 12229
rect 13193 12189 13205 12223
rect 13239 12220 13251 12223
rect 13354 12220 13360 12232
rect 13239 12192 13360 12220
rect 13239 12189 13251 12192
rect 13193 12183 13251 12189
rect 9214 12152 9220 12164
rect 8864 12124 9220 12152
rect 9214 12112 9220 12124
rect 9272 12112 9278 12164
rect 11348 12152 11376 12183
rect 13354 12180 13360 12192
rect 13412 12180 13418 12232
rect 13556 12229 13584 12384
rect 18138 12316 18144 12368
rect 18196 12356 18202 12368
rect 18877 12359 18935 12365
rect 18877 12356 18889 12359
rect 18196 12328 18889 12356
rect 18196 12316 18202 12328
rect 18877 12325 18889 12328
rect 18923 12325 18935 12359
rect 18877 12319 18935 12325
rect 17494 12288 17500 12300
rect 15396 12260 17500 12288
rect 13541 12223 13599 12229
rect 13541 12189 13553 12223
rect 13587 12220 13599 12223
rect 15217 12223 15275 12229
rect 13587 12192 13676 12220
rect 13587 12189 13599 12192
rect 13541 12183 13599 12189
rect 9646 12124 11376 12152
rect 5721 12087 5779 12093
rect 5721 12084 5733 12087
rect 2056 12056 5733 12084
rect 5721 12053 5733 12056
rect 5767 12053 5779 12087
rect 5721 12047 5779 12053
rect 5905 12087 5963 12093
rect 5905 12053 5917 12087
rect 5951 12084 5963 12087
rect 6270 12084 6276 12096
rect 5951 12056 6276 12084
rect 5951 12053 5963 12056
rect 5905 12047 5963 12053
rect 6270 12044 6276 12056
rect 6328 12044 6334 12096
rect 7377 12087 7435 12093
rect 7377 12053 7389 12087
rect 7423 12084 7435 12087
rect 7466 12084 7472 12096
rect 7423 12056 7472 12084
rect 7423 12053 7435 12056
rect 7377 12047 7435 12053
rect 7466 12044 7472 12056
rect 7524 12084 7530 12096
rect 9646 12084 9674 12124
rect 11882 12112 11888 12164
rect 11940 12152 11946 12164
rect 11977 12155 12035 12161
rect 11977 12152 11989 12155
rect 11940 12124 11989 12152
rect 11940 12112 11946 12124
rect 11977 12121 11989 12124
rect 12023 12121 12035 12155
rect 11977 12115 12035 12121
rect 13648 12096 13676 12192
rect 15217 12189 15229 12223
rect 15263 12220 15275 12223
rect 15396 12220 15424 12260
rect 17494 12248 17500 12260
rect 17552 12248 17558 12300
rect 17586 12248 17592 12300
rect 17644 12288 17650 12300
rect 17644 12260 18828 12288
rect 17644 12248 17650 12260
rect 15263 12192 15424 12220
rect 15473 12223 15531 12229
rect 15263 12189 15275 12192
rect 15217 12183 15275 12189
rect 15473 12189 15485 12223
rect 15519 12220 15531 12223
rect 15657 12223 15715 12229
rect 15657 12220 15669 12223
rect 15519 12192 15669 12220
rect 15519 12189 15531 12192
rect 15473 12183 15531 12189
rect 15657 12189 15669 12192
rect 15703 12189 15715 12223
rect 15657 12183 15715 12189
rect 15749 12223 15807 12229
rect 15749 12189 15761 12223
rect 15795 12189 15807 12223
rect 15749 12183 15807 12189
rect 7524 12056 9674 12084
rect 7524 12044 7530 12056
rect 10226 12044 10232 12096
rect 10284 12044 10290 12096
rect 11330 12044 11336 12096
rect 11388 12084 11394 12096
rect 11517 12087 11575 12093
rect 11517 12084 11529 12087
rect 11388 12056 11529 12084
rect 11388 12044 11394 12056
rect 11517 12053 11529 12056
rect 11563 12053 11575 12087
rect 11517 12047 11575 12053
rect 13630 12044 13636 12096
rect 13688 12044 13694 12096
rect 14093 12087 14151 12093
rect 14093 12053 14105 12087
rect 14139 12084 14151 12087
rect 14366 12084 14372 12096
rect 14139 12056 14372 12084
rect 14139 12053 14151 12056
rect 14093 12047 14151 12053
rect 14366 12044 14372 12056
rect 14424 12044 14430 12096
rect 15764 12084 15792 12183
rect 16022 12180 16028 12232
rect 16080 12180 16086 12232
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12220 18015 12223
rect 18138 12220 18144 12232
rect 18003 12192 18144 12220
rect 18003 12189 18015 12192
rect 17957 12183 18015 12189
rect 18138 12180 18144 12192
rect 18196 12180 18202 12232
rect 18800 12229 18828 12260
rect 18509 12223 18567 12229
rect 18509 12189 18521 12223
rect 18555 12220 18567 12223
rect 18785 12223 18843 12229
rect 18555 12192 18736 12220
rect 18555 12189 18567 12192
rect 18509 12183 18567 12189
rect 16666 12112 16672 12164
rect 16724 12152 16730 12164
rect 18708 12152 18736 12192
rect 18785 12189 18797 12223
rect 18831 12189 18843 12223
rect 18785 12183 18843 12189
rect 19058 12180 19064 12232
rect 19116 12180 19122 12232
rect 19260 12229 19288 12396
rect 22649 12393 22661 12427
rect 22695 12424 22707 12427
rect 23106 12424 23112 12436
rect 22695 12396 23112 12424
rect 22695 12393 22707 12396
rect 22649 12387 22707 12393
rect 23106 12384 23112 12396
rect 23164 12424 23170 12436
rect 23382 12424 23388 12436
rect 23164 12396 23388 12424
rect 23164 12384 23170 12396
rect 23382 12384 23388 12396
rect 23440 12384 23446 12436
rect 21174 12248 21180 12300
rect 21232 12288 21238 12300
rect 21818 12288 21824 12300
rect 21232 12260 21824 12288
rect 21232 12248 21238 12260
rect 21818 12248 21824 12260
rect 21876 12248 21882 12300
rect 19245 12223 19303 12229
rect 19245 12189 19257 12223
rect 19291 12189 19303 12223
rect 19245 12183 19303 12189
rect 19702 12180 19708 12232
rect 19760 12220 19766 12232
rect 23474 12220 23480 12232
rect 19760 12192 23480 12220
rect 19760 12180 19766 12192
rect 23474 12180 23480 12192
rect 23532 12180 23538 12232
rect 20438 12152 20444 12164
rect 16724 12124 18644 12152
rect 18708 12124 20444 12152
rect 16724 12112 16730 12124
rect 16114 12084 16120 12096
rect 15764 12056 16120 12084
rect 16114 12044 16120 12056
rect 16172 12084 16178 12096
rect 17313 12087 17371 12093
rect 17313 12084 17325 12087
rect 16172 12056 17325 12084
rect 16172 12044 16178 12056
rect 17313 12053 17325 12056
rect 17359 12084 17371 12087
rect 18414 12084 18420 12096
rect 17359 12056 18420 12084
rect 17359 12053 17371 12056
rect 17313 12047 17371 12053
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 18616 12093 18644 12124
rect 20438 12112 20444 12124
rect 20496 12112 20502 12164
rect 21177 12155 21235 12161
rect 21177 12152 21189 12155
rect 20548 12124 21189 12152
rect 20548 12096 20576 12124
rect 21177 12121 21189 12124
rect 21223 12121 21235 12155
rect 21177 12115 21235 12121
rect 22066 12124 22876 12152
rect 18601 12087 18659 12093
rect 18601 12053 18613 12087
rect 18647 12053 18659 12087
rect 18601 12047 18659 12053
rect 20530 12044 20536 12096
rect 20588 12044 20594 12096
rect 21082 12044 21088 12096
rect 21140 12084 21146 12096
rect 22066 12084 22094 12124
rect 22848 12096 22876 12124
rect 21140 12056 22094 12084
rect 21140 12044 21146 12056
rect 22830 12044 22836 12096
rect 22888 12044 22894 12096
rect 1104 11994 23828 12016
rect 1104 11942 2658 11994
rect 2710 11942 2722 11994
rect 2774 11942 2786 11994
rect 2838 11942 2850 11994
rect 2902 11942 2914 11994
rect 2966 11942 2978 11994
rect 3030 11942 8658 11994
rect 8710 11942 8722 11994
rect 8774 11942 8786 11994
rect 8838 11942 8850 11994
rect 8902 11942 8914 11994
rect 8966 11942 8978 11994
rect 9030 11942 14658 11994
rect 14710 11942 14722 11994
rect 14774 11942 14786 11994
rect 14838 11942 14850 11994
rect 14902 11942 14914 11994
rect 14966 11942 14978 11994
rect 15030 11942 20658 11994
rect 20710 11942 20722 11994
rect 20774 11942 20786 11994
rect 20838 11942 20850 11994
rect 20902 11942 20914 11994
rect 20966 11942 20978 11994
rect 21030 11942 23828 11994
rect 1104 11920 23828 11942
rect 1578 11840 1584 11892
rect 1636 11840 1642 11892
rect 11054 11840 11060 11892
rect 11112 11880 11118 11892
rect 11149 11883 11207 11889
rect 11149 11880 11161 11883
rect 11112 11852 11161 11880
rect 11112 11840 11118 11852
rect 11149 11849 11161 11852
rect 11195 11849 11207 11883
rect 15746 11880 15752 11892
rect 11149 11843 11207 11849
rect 11348 11852 15752 11880
rect 1596 11753 1624 11840
rect 1762 11772 1768 11824
rect 1820 11812 1826 11824
rect 2102 11815 2160 11821
rect 2102 11812 2114 11815
rect 1820 11784 2114 11812
rect 1820 11772 1826 11784
rect 2102 11781 2114 11784
rect 2148 11781 2160 11815
rect 2102 11775 2160 11781
rect 2498 11772 2504 11824
rect 2556 11812 2562 11824
rect 7837 11815 7895 11821
rect 7837 11812 7849 11815
rect 2556 11784 7849 11812
rect 2556 11772 2562 11784
rect 7837 11781 7849 11784
rect 7883 11781 7895 11815
rect 7837 11775 7895 11781
rect 9766 11772 9772 11824
rect 9824 11812 9830 11824
rect 9922 11815 9980 11821
rect 9922 11812 9934 11815
rect 9824 11784 9934 11812
rect 9824 11772 9830 11784
rect 9922 11781 9934 11784
rect 9968 11781 9980 11815
rect 9922 11775 9980 11781
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 3234 11704 3240 11756
rect 3292 11744 3298 11756
rect 3585 11747 3643 11753
rect 3585 11744 3597 11747
rect 3292 11716 3597 11744
rect 3292 11704 3298 11716
rect 3585 11713 3597 11716
rect 3631 11713 3643 11747
rect 3585 11707 3643 11713
rect 5902 11704 5908 11756
rect 5960 11753 5966 11756
rect 5960 11747 5983 11753
rect 5971 11713 5983 11747
rect 5960 11707 5983 11713
rect 5960 11704 5966 11707
rect 6086 11704 6092 11756
rect 6144 11744 6150 11756
rect 6181 11747 6239 11753
rect 6181 11744 6193 11747
rect 6144 11716 6193 11744
rect 6144 11704 6150 11716
rect 6181 11713 6193 11716
rect 6227 11713 6239 11747
rect 6181 11707 6239 11713
rect 6632 11747 6690 11753
rect 6632 11713 6644 11747
rect 6678 11744 6690 11747
rect 6678 11716 9628 11744
rect 6678 11713 6690 11716
rect 6632 11707 6690 11713
rect 1486 11636 1492 11688
rect 1544 11676 1550 11688
rect 1857 11679 1915 11685
rect 1857 11676 1869 11679
rect 1544 11648 1869 11676
rect 1544 11636 1550 11648
rect 1857 11645 1869 11648
rect 1903 11645 1915 11679
rect 1857 11639 1915 11645
rect 3050 11636 3056 11688
rect 3108 11676 3114 11688
rect 3329 11679 3387 11685
rect 3329 11676 3341 11679
rect 3108 11648 3341 11676
rect 3108 11636 3114 11648
rect 3329 11645 3341 11648
rect 3375 11645 3387 11679
rect 3329 11639 3387 11645
rect 6362 11636 6368 11688
rect 6420 11636 6426 11688
rect 9600 11676 9628 11716
rect 9674 11704 9680 11756
rect 9732 11704 9738 11756
rect 10502 11744 10508 11756
rect 9784 11716 10508 11744
rect 9784 11676 9812 11716
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 11348 11753 11376 11852
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 21082 11880 21088 11892
rect 18340 11852 21088 11880
rect 12802 11772 12808 11824
rect 12860 11812 12866 11824
rect 13081 11815 13139 11821
rect 13081 11812 13093 11815
rect 12860 11784 13093 11812
rect 12860 11772 12866 11784
rect 13081 11781 13093 11784
rect 13127 11781 13139 11815
rect 13081 11775 13139 11781
rect 14829 11815 14887 11821
rect 14829 11781 14841 11815
rect 14875 11812 14887 11815
rect 15102 11812 15108 11824
rect 14875 11784 15108 11812
rect 14875 11781 14887 11784
rect 14829 11775 14887 11781
rect 15102 11772 15108 11784
rect 15160 11772 15166 11824
rect 11333 11747 11391 11753
rect 11333 11713 11345 11747
rect 11379 11713 11391 11747
rect 11333 11707 11391 11713
rect 11606 11704 11612 11756
rect 11664 11704 11670 11756
rect 11698 11704 11704 11756
rect 11756 11744 11762 11756
rect 11865 11747 11923 11753
rect 11865 11744 11877 11747
rect 11756 11716 11877 11744
rect 11756 11704 11762 11716
rect 11865 11713 11877 11716
rect 11911 11713 11923 11747
rect 11865 11707 11923 11713
rect 15188 11747 15246 11753
rect 15188 11713 15200 11747
rect 15234 11744 15246 11747
rect 15562 11744 15568 11756
rect 15234 11716 15568 11744
rect 15234 11713 15246 11716
rect 15188 11707 15246 11713
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 18340 11744 18368 11852
rect 21082 11840 21088 11852
rect 21140 11840 21146 11892
rect 21542 11840 21548 11892
rect 21600 11840 21606 11892
rect 21634 11840 21640 11892
rect 21692 11880 21698 11892
rect 23385 11883 23443 11889
rect 23385 11880 23397 11883
rect 21692 11852 23397 11880
rect 21692 11840 21698 11852
rect 23385 11849 23397 11852
rect 23431 11849 23443 11883
rect 23385 11843 23443 11849
rect 18417 11815 18475 11821
rect 18417 11781 18429 11815
rect 18463 11812 18475 11815
rect 20530 11812 20536 11824
rect 18463 11784 20536 11812
rect 18463 11781 18475 11784
rect 18417 11775 18475 11781
rect 20530 11772 20536 11784
rect 20588 11772 20594 11824
rect 21358 11772 21364 11824
rect 21416 11812 21422 11824
rect 22088 11815 22146 11821
rect 21416 11784 21680 11812
rect 21416 11772 21422 11784
rect 21652 11756 21680 11784
rect 22088 11781 22100 11815
rect 22134 11812 22146 11815
rect 22554 11812 22560 11824
rect 22134 11784 22560 11812
rect 22134 11781 22146 11784
rect 22088 11775 22146 11781
rect 22554 11772 22560 11784
rect 22612 11772 22618 11824
rect 18509 11747 18567 11753
rect 18509 11744 18521 11747
rect 18340 11716 18521 11744
rect 18509 11713 18521 11716
rect 18555 11713 18567 11747
rect 18509 11707 18567 11713
rect 18598 11704 18604 11756
rect 18656 11744 18662 11756
rect 18765 11747 18823 11753
rect 18765 11744 18777 11747
rect 18656 11716 18777 11744
rect 18656 11704 18662 11716
rect 18765 11713 18777 11716
rect 18811 11713 18823 11747
rect 18765 11707 18823 11713
rect 21105 11747 21163 11753
rect 21105 11713 21117 11747
rect 21151 11744 21163 11747
rect 21151 11716 21588 11744
rect 21151 11713 21163 11716
rect 21105 11707 21163 11713
rect 11238 11676 11244 11688
rect 9600 11648 9812 11676
rect 11072 11648 11244 11676
rect 1762 11568 1768 11620
rect 1820 11568 1826 11620
rect 4338 11568 4344 11620
rect 4396 11608 4402 11620
rect 11072 11617 11100 11648
rect 11238 11636 11244 11648
rect 11296 11636 11302 11688
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 21361 11679 21419 11685
rect 21361 11645 21373 11679
rect 21407 11645 21419 11679
rect 21560 11676 21588 11716
rect 21634 11704 21640 11756
rect 21692 11704 21698 11756
rect 21910 11744 21916 11756
rect 21744 11716 21916 11744
rect 21744 11676 21772 11716
rect 21910 11704 21916 11716
rect 21968 11704 21974 11756
rect 23290 11704 23296 11756
rect 23348 11704 23354 11756
rect 21560 11648 21772 11676
rect 21361 11639 21419 11645
rect 4801 11611 4859 11617
rect 4801 11608 4813 11611
rect 4396 11580 4813 11608
rect 4396 11568 4402 11580
rect 4801 11577 4813 11580
rect 4847 11577 4859 11611
rect 4801 11571 4859 11577
rect 11057 11611 11115 11617
rect 11057 11577 11069 11611
rect 11103 11577 11115 11611
rect 11057 11571 11115 11577
rect 3237 11543 3295 11549
rect 3237 11509 3249 11543
rect 3283 11540 3295 11543
rect 3326 11540 3332 11552
rect 3283 11512 3332 11540
rect 3283 11509 3295 11512
rect 3237 11503 3295 11509
rect 3326 11500 3332 11512
rect 3384 11500 3390 11552
rect 3510 11500 3516 11552
rect 3568 11540 3574 11552
rect 4709 11543 4767 11549
rect 4709 11540 4721 11543
rect 3568 11512 4721 11540
rect 3568 11500 3574 11512
rect 4709 11509 4721 11512
rect 4755 11509 4767 11543
rect 4709 11503 4767 11509
rect 7650 11500 7656 11552
rect 7708 11540 7714 11552
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 7708 11512 7757 11540
rect 7708 11500 7714 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 7745 11503 7803 11509
rect 8478 11500 8484 11552
rect 8536 11540 8542 11552
rect 9122 11540 9128 11552
rect 8536 11512 9128 11540
rect 8536 11500 8542 11512
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 11146 11500 11152 11552
rect 11204 11540 11210 11552
rect 11790 11540 11796 11552
rect 11204 11512 11796 11540
rect 11204 11500 11210 11512
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 12986 11500 12992 11552
rect 13044 11500 13050 11552
rect 14936 11540 14964 11639
rect 16301 11611 16359 11617
rect 16301 11577 16313 11611
rect 16347 11608 16359 11611
rect 17586 11608 17592 11620
rect 16347 11580 17592 11608
rect 16347 11577 16359 11580
rect 16301 11571 16359 11577
rect 17586 11568 17592 11580
rect 17644 11568 17650 11620
rect 16206 11540 16212 11552
rect 14936 11512 16212 11540
rect 16206 11500 16212 11512
rect 16264 11500 16270 11552
rect 16758 11500 16764 11552
rect 16816 11540 16822 11552
rect 16945 11543 17003 11549
rect 16945 11540 16957 11543
rect 16816 11512 16957 11540
rect 16816 11500 16822 11512
rect 16945 11509 16957 11512
rect 16991 11509 17003 11543
rect 16945 11503 17003 11509
rect 19794 11500 19800 11552
rect 19852 11540 19858 11552
rect 19889 11543 19947 11549
rect 19889 11540 19901 11543
rect 19852 11512 19901 11540
rect 19852 11500 19858 11512
rect 19889 11509 19901 11512
rect 19935 11509 19947 11543
rect 19889 11503 19947 11509
rect 19981 11543 20039 11549
rect 19981 11509 19993 11543
rect 20027 11540 20039 11543
rect 21174 11540 21180 11552
rect 20027 11512 21180 11540
rect 20027 11509 20039 11512
rect 19981 11503 20039 11509
rect 21174 11500 21180 11512
rect 21232 11500 21238 11552
rect 21376 11540 21404 11639
rect 21818 11636 21824 11688
rect 21876 11636 21882 11688
rect 23014 11568 23020 11620
rect 23072 11608 23078 11620
rect 23201 11611 23259 11617
rect 23201 11608 23213 11611
rect 23072 11580 23213 11608
rect 23072 11568 23078 11580
rect 23201 11577 23213 11580
rect 23247 11577 23259 11611
rect 23201 11571 23259 11577
rect 22462 11540 22468 11552
rect 21376 11512 22468 11540
rect 22462 11500 22468 11512
rect 22520 11500 22526 11552
rect 1104 11450 23828 11472
rect 1104 11398 1918 11450
rect 1970 11398 1982 11450
rect 2034 11398 2046 11450
rect 2098 11398 2110 11450
rect 2162 11398 2174 11450
rect 2226 11398 2238 11450
rect 2290 11398 7918 11450
rect 7970 11398 7982 11450
rect 8034 11398 8046 11450
rect 8098 11398 8110 11450
rect 8162 11398 8174 11450
rect 8226 11398 8238 11450
rect 8290 11398 13918 11450
rect 13970 11398 13982 11450
rect 14034 11398 14046 11450
rect 14098 11398 14110 11450
rect 14162 11398 14174 11450
rect 14226 11398 14238 11450
rect 14290 11398 19918 11450
rect 19970 11398 19982 11450
rect 20034 11398 20046 11450
rect 20098 11398 20110 11450
rect 20162 11398 20174 11450
rect 20226 11398 20238 11450
rect 20290 11398 23828 11450
rect 1104 11376 23828 11398
rect 2133 11339 2191 11345
rect 2133 11305 2145 11339
rect 2179 11336 2191 11339
rect 2179 11308 5396 11336
rect 2179 11305 2191 11308
rect 2133 11299 2191 11305
rect 5368 11268 5396 11308
rect 5626 11296 5632 11348
rect 5684 11336 5690 11348
rect 5813 11339 5871 11345
rect 5813 11336 5825 11339
rect 5684 11308 5825 11336
rect 5684 11296 5690 11308
rect 5813 11305 5825 11308
rect 5859 11305 5871 11339
rect 5813 11299 5871 11305
rect 8757 11339 8815 11345
rect 8757 11305 8769 11339
rect 8803 11336 8815 11339
rect 11698 11336 11704 11348
rect 8803 11308 11704 11336
rect 8803 11305 8815 11308
rect 8757 11299 8815 11305
rect 11698 11296 11704 11308
rect 11756 11296 11762 11348
rect 12161 11339 12219 11345
rect 12161 11305 12173 11339
rect 12207 11336 12219 11339
rect 12802 11336 12808 11348
rect 12207 11308 12808 11336
rect 12207 11305 12219 11308
rect 12161 11299 12219 11305
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 13262 11296 13268 11348
rect 13320 11336 13326 11348
rect 13817 11339 13875 11345
rect 13320 11308 13768 11336
rect 13320 11296 13326 11308
rect 11241 11271 11299 11277
rect 5368 11240 5856 11268
rect 5828 11212 5856 11240
rect 11241 11237 11253 11271
rect 11287 11268 11299 11271
rect 11606 11268 11612 11280
rect 11287 11240 11612 11268
rect 11287 11237 11299 11240
rect 11241 11231 11299 11237
rect 11606 11228 11612 11240
rect 11664 11228 11670 11280
rect 13740 11268 13768 11308
rect 13817 11305 13829 11339
rect 13863 11336 13875 11339
rect 15470 11336 15476 11348
rect 13863 11308 15476 11336
rect 13863 11305 13875 11308
rect 13817 11299 13875 11305
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 23290 11336 23296 11348
rect 16684 11308 23296 11336
rect 13740 11240 14688 11268
rect 3326 11160 3332 11212
rect 3384 11200 3390 11212
rect 3602 11200 3608 11212
rect 3384 11172 3608 11200
rect 3384 11160 3390 11172
rect 3602 11160 3608 11172
rect 3660 11160 3666 11212
rect 4080 11172 4568 11200
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11101 1639 11135
rect 1581 11095 1639 11101
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11132 2283 11135
rect 2314 11132 2320 11144
rect 2271 11104 2320 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 1596 11064 1624 11095
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 4080 11132 4108 11172
rect 2424 11104 4108 11132
rect 2424 11064 2452 11104
rect 4430 11092 4436 11144
rect 4488 11092 4494 11144
rect 4540 11132 4568 11172
rect 5810 11160 5816 11212
rect 5868 11160 5874 11212
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11200 11391 11203
rect 11977 11203 12035 11209
rect 11977 11200 11989 11203
rect 11379 11172 11989 11200
rect 11379 11169 11391 11172
rect 11333 11163 11391 11169
rect 11977 11169 11989 11172
rect 12023 11169 12035 11203
rect 11977 11163 12035 11169
rect 13541 11203 13599 11209
rect 13541 11169 13553 11203
rect 13587 11200 13599 11203
rect 14090 11200 14096 11212
rect 13587 11172 14096 11200
rect 13587 11169 13599 11172
rect 13541 11163 13599 11169
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 14660 11209 14688 11240
rect 15286 11228 15292 11280
rect 15344 11268 15350 11280
rect 16684 11268 16712 11308
rect 23290 11296 23296 11308
rect 23348 11296 23354 11348
rect 15344 11240 16712 11268
rect 16761 11271 16819 11277
rect 15344 11228 15350 11240
rect 16761 11237 16773 11271
rect 16807 11237 16819 11271
rect 16761 11231 16819 11237
rect 19613 11271 19671 11277
rect 19613 11237 19625 11271
rect 19659 11268 19671 11271
rect 19659 11240 20300 11268
rect 19659 11237 19671 11240
rect 19613 11231 19671 11237
rect 14645 11203 14703 11209
rect 14645 11169 14657 11203
rect 14691 11169 14703 11203
rect 14645 11163 14703 11169
rect 16666 11160 16672 11212
rect 16724 11200 16730 11212
rect 16776 11200 16804 11231
rect 16724 11172 16804 11200
rect 16724 11160 16730 11172
rect 17126 11160 17132 11212
rect 17184 11200 17190 11212
rect 18506 11200 18512 11212
rect 17184 11172 18512 11200
rect 17184 11160 17190 11172
rect 18506 11160 18512 11172
rect 18564 11200 18570 11212
rect 19245 11203 19303 11209
rect 19245 11200 19257 11203
rect 18564 11172 19257 11200
rect 18564 11160 18570 11172
rect 19245 11169 19257 11172
rect 19291 11169 19303 11203
rect 19245 11163 19303 11169
rect 19702 11160 19708 11212
rect 19760 11160 19766 11212
rect 5442 11132 5448 11144
rect 4540 11104 5448 11132
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 5534 11092 5540 11144
rect 5592 11132 5598 11144
rect 6089 11135 6147 11141
rect 6089 11132 6101 11135
rect 5592 11104 6101 11132
rect 5592 11092 5598 11104
rect 6089 11101 6101 11104
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 7374 11092 7380 11144
rect 7432 11092 7438 11144
rect 7650 11141 7656 11144
rect 7644 11132 7656 11141
rect 7611 11104 7656 11132
rect 7644 11095 7656 11104
rect 7650 11092 7656 11095
rect 7708 11092 7714 11144
rect 10778 11092 10784 11144
rect 10836 11132 10842 11144
rect 11425 11135 11483 11141
rect 11425 11132 11437 11135
rect 10836 11104 11437 11132
rect 10836 11092 10842 11104
rect 11425 11101 11437 11104
rect 11471 11101 11483 11135
rect 11425 11095 11483 11101
rect 12986 11092 12992 11144
rect 13044 11132 13050 11144
rect 13262 11132 13268 11144
rect 13320 11141 13326 11144
rect 13044 11104 13268 11132
rect 13044 11092 13050 11104
rect 13262 11092 13268 11104
rect 13320 11095 13332 11141
rect 13320 11092 13326 11095
rect 13630 11092 13636 11144
rect 13688 11128 13694 11144
rect 15102 11132 15108 11144
rect 13740 11128 15108 11132
rect 13688 11104 15108 11128
rect 13688 11100 13768 11104
rect 13688 11092 13694 11100
rect 1596 11036 2452 11064
rect 2492 11067 2550 11073
rect 2492 11033 2504 11067
rect 2538 11064 2550 11067
rect 3234 11064 3240 11076
rect 2538 11036 3240 11064
rect 2538 11033 2550 11036
rect 2492 11027 2550 11033
rect 3234 11024 3240 11036
rect 3292 11024 3298 11076
rect 3694 11064 3700 11076
rect 3620 11036 3700 11064
rect 3620 11005 3648 11036
rect 3694 11024 3700 11036
rect 3752 11024 3758 11076
rect 4522 11024 4528 11076
rect 4580 11064 4586 11076
rect 4678 11067 4736 11073
rect 4678 11064 4690 11067
rect 4580 11036 4690 11064
rect 4580 11024 4586 11036
rect 4678 11033 4690 11036
rect 4724 11033 4736 11067
rect 4678 11027 4736 11033
rect 4798 11024 4804 11076
rect 4856 11064 4862 11076
rect 6457 11067 6515 11073
rect 6457 11064 6469 11067
rect 4856 11036 6469 11064
rect 4856 11024 4862 11036
rect 6457 11033 6469 11036
rect 6503 11033 6515 11067
rect 6457 11027 6515 11033
rect 8941 11067 8999 11073
rect 8941 11033 8953 11067
rect 8987 11064 8999 11067
rect 9122 11064 9128 11076
rect 8987 11036 9128 11064
rect 8987 11033 8999 11036
rect 8941 11027 8999 11033
rect 9122 11024 9128 11036
rect 9180 11024 9186 11076
rect 9214 11024 9220 11076
rect 9272 11064 9278 11076
rect 10505 11067 10563 11073
rect 10505 11064 10517 11067
rect 9272 11036 10517 11064
rect 9272 11024 9278 11036
rect 10505 11033 10517 11036
rect 10551 11033 10563 11067
rect 10505 11027 10563 11033
rect 10873 11067 10931 11073
rect 10873 11033 10885 11067
rect 10919 11064 10931 11067
rect 11146 11064 11152 11076
rect 10919 11036 11152 11064
rect 10919 11033 10931 11036
rect 10873 11027 10931 11033
rect 11146 11024 11152 11036
rect 11204 11024 11210 11076
rect 11256 11036 11560 11064
rect 3605 10999 3663 11005
rect 3605 10965 3617 10999
rect 3651 10965 3663 10999
rect 3605 10959 3663 10965
rect 7466 10956 7472 11008
rect 7524 10996 7530 11008
rect 11256 10996 11284 11036
rect 7524 10968 11284 10996
rect 11532 10996 11560 11036
rect 12084 11036 12296 11064
rect 12084 10996 12112 11036
rect 11532 10968 12112 10996
rect 12268 10996 12296 11036
rect 13740 10996 13768 11100
rect 15102 11092 15108 11104
rect 15160 11092 15166 11144
rect 16577 11135 16635 11141
rect 16577 11101 16589 11135
rect 16623 11132 16635 11135
rect 18877 11135 18935 11141
rect 18877 11132 18889 11135
rect 16623 11104 18889 11132
rect 16623 11101 16635 11104
rect 16577 11095 16635 11101
rect 18877 11101 18889 11104
rect 18923 11132 18935 11135
rect 19797 11135 19855 11141
rect 19797 11132 19809 11135
rect 18923 11104 19809 11132
rect 18923 11101 18935 11104
rect 18877 11095 18935 11101
rect 19797 11101 19809 11104
rect 19843 11101 19855 11135
rect 19797 11095 19855 11101
rect 14093 11067 14151 11073
rect 14093 11033 14105 11067
rect 14139 11064 14151 11067
rect 14274 11064 14280 11076
rect 14139 11036 14280 11064
rect 14139 11033 14151 11036
rect 14093 11027 14151 11033
rect 14274 11024 14280 11036
rect 14332 11024 14338 11076
rect 15378 11024 15384 11076
rect 15436 11064 15442 11076
rect 17313 11067 17371 11073
rect 17313 11064 17325 11067
rect 15436 11036 17080 11064
rect 15436 11024 15442 11036
rect 12268 10968 13768 10996
rect 16669 10999 16727 11005
rect 7524 10956 7530 10968
rect 16669 10965 16681 10999
rect 16715 10996 16727 10999
rect 16942 10996 16948 11008
rect 16715 10968 16948 10996
rect 16715 10965 16727 10968
rect 16669 10959 16727 10965
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 17052 10996 17080 11036
rect 17236 11036 17325 11064
rect 17236 10996 17264 11036
rect 17313 11033 17325 11036
rect 17359 11033 17371 11067
rect 20272 11064 20300 11240
rect 22002 11228 22008 11280
rect 22060 11228 22066 11280
rect 21542 11160 21548 11212
rect 21600 11200 21606 11212
rect 22020 11200 22048 11228
rect 21600 11172 22048 11200
rect 21600 11160 21606 11172
rect 20346 11092 20352 11144
rect 20404 11132 20410 11144
rect 20404 11104 22876 11132
rect 20404 11092 20410 11104
rect 22094 11064 22100 11076
rect 20272 11036 22100 11064
rect 17313 11027 17371 11033
rect 22094 11024 22100 11036
rect 22152 11024 22158 11076
rect 22750 11067 22808 11073
rect 22750 11064 22762 11067
rect 22204 11036 22762 11064
rect 17052 10968 17264 10996
rect 17770 10956 17776 11008
rect 17828 10996 17834 11008
rect 19610 10996 19616 11008
rect 17828 10968 19616 10996
rect 17828 10956 17834 10968
rect 19610 10956 19616 10968
rect 19668 10956 19674 11008
rect 21450 10956 21456 11008
rect 21508 10996 21514 11008
rect 21637 10999 21695 11005
rect 21637 10996 21649 10999
rect 21508 10968 21649 10996
rect 21508 10956 21514 10968
rect 21637 10965 21649 10968
rect 21683 10965 21695 10999
rect 21637 10959 21695 10965
rect 22002 10956 22008 11008
rect 22060 10996 22066 11008
rect 22204 10996 22232 11036
rect 22750 11033 22762 11036
rect 22796 11033 22808 11067
rect 22848 11064 22876 11104
rect 23014 11092 23020 11144
rect 23072 11092 23078 11144
rect 23106 11092 23112 11144
rect 23164 11092 23170 11144
rect 23201 11135 23259 11141
rect 23201 11101 23213 11135
rect 23247 11101 23259 11135
rect 23201 11095 23259 11101
rect 23216 11064 23244 11095
rect 22848 11036 23244 11064
rect 22750 11027 22808 11033
rect 22060 10968 22232 10996
rect 22060 10956 22066 10968
rect 1104 10906 23828 10928
rect 1104 10854 2658 10906
rect 2710 10854 2722 10906
rect 2774 10854 2786 10906
rect 2838 10854 2850 10906
rect 2902 10854 2914 10906
rect 2966 10854 2978 10906
rect 3030 10854 8658 10906
rect 8710 10854 8722 10906
rect 8774 10854 8786 10906
rect 8838 10854 8850 10906
rect 8902 10854 8914 10906
rect 8966 10854 8978 10906
rect 9030 10854 14658 10906
rect 14710 10854 14722 10906
rect 14774 10854 14786 10906
rect 14838 10854 14850 10906
rect 14902 10854 14914 10906
rect 14966 10854 14978 10906
rect 15030 10854 20658 10906
rect 20710 10854 20722 10906
rect 20774 10854 20786 10906
rect 20838 10854 20850 10906
rect 20902 10854 20914 10906
rect 20966 10854 20978 10906
rect 21030 10854 23828 10906
rect 1104 10832 23828 10854
rect 4617 10795 4675 10801
rect 1780 10764 3536 10792
rect 1210 10616 1216 10668
rect 1268 10616 1274 10668
rect 1489 10659 1547 10665
rect 1489 10625 1501 10659
rect 1535 10656 1547 10659
rect 1780 10656 1808 10764
rect 2222 10684 2228 10736
rect 2280 10724 2286 10736
rect 2498 10724 2504 10736
rect 2280 10696 2504 10724
rect 2280 10684 2286 10696
rect 2498 10684 2504 10696
rect 2556 10684 2562 10736
rect 3508 10724 3536 10764
rect 4617 10761 4629 10795
rect 4663 10792 4675 10795
rect 5534 10792 5540 10804
rect 4663 10764 5540 10792
rect 4663 10761 4675 10764
rect 4617 10755 4675 10761
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 13814 10792 13820 10804
rect 11164 10764 13820 10792
rect 7282 10724 7288 10736
rect 2746 10696 3464 10724
rect 3508 10696 7288 10724
rect 1535 10628 1808 10656
rect 1535 10625 1547 10628
rect 1489 10619 1547 10625
rect 1854 10616 1860 10668
rect 1912 10656 1918 10668
rect 2021 10659 2079 10665
rect 2021 10656 2033 10659
rect 1912 10628 2033 10656
rect 1912 10616 1918 10628
rect 2021 10625 2033 10628
rect 2067 10625 2079 10659
rect 2021 10619 2079 10625
rect 2590 10616 2596 10668
rect 2648 10656 2654 10668
rect 2746 10656 2774 10696
rect 2648 10628 2774 10656
rect 2648 10616 2654 10628
rect 3142 10616 3148 10668
rect 3200 10616 3206 10668
rect 3237 10659 3295 10665
rect 3237 10625 3249 10659
rect 3283 10656 3295 10659
rect 3326 10656 3332 10668
rect 3283 10628 3332 10656
rect 3283 10625 3295 10628
rect 3237 10619 3295 10625
rect 3326 10616 3332 10628
rect 3384 10616 3390 10668
rect 3436 10656 3464 10696
rect 7282 10684 7288 10696
rect 7340 10684 7346 10736
rect 7466 10684 7472 10736
rect 7524 10684 7530 10736
rect 8478 10684 8484 10736
rect 8536 10684 8542 10736
rect 3493 10659 3551 10665
rect 3493 10656 3505 10659
rect 3436 10628 3505 10656
rect 3493 10625 3505 10628
rect 3539 10625 3551 10659
rect 3493 10619 3551 10625
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 5057 10659 5115 10665
rect 5057 10656 5069 10659
rect 3936 10628 5069 10656
rect 3936 10616 3942 10628
rect 5057 10625 5069 10628
rect 5103 10625 5115 10659
rect 5057 10619 5115 10625
rect 6454 10616 6460 10668
rect 6512 10656 6518 10668
rect 7484 10656 7512 10684
rect 6512 10628 7512 10656
rect 6512 10616 6518 10628
rect 7834 10616 7840 10668
rect 7892 10656 7898 10668
rect 11164 10665 11192 10764
rect 13814 10752 13820 10764
rect 13872 10752 13878 10804
rect 15473 10795 15531 10801
rect 15473 10761 15485 10795
rect 15519 10792 15531 10795
rect 15562 10792 15568 10804
rect 15519 10764 15568 10792
rect 15519 10761 15531 10764
rect 15473 10755 15531 10761
rect 15562 10752 15568 10764
rect 15620 10752 15626 10804
rect 16209 10795 16267 10801
rect 16209 10761 16221 10795
rect 16255 10792 16267 10795
rect 16574 10792 16580 10804
rect 16255 10764 16580 10792
rect 16255 10761 16267 10764
rect 16209 10755 16267 10761
rect 16574 10752 16580 10764
rect 16632 10752 16638 10804
rect 16761 10795 16819 10801
rect 16761 10761 16773 10795
rect 16807 10792 16819 10795
rect 17310 10792 17316 10804
rect 16807 10764 17316 10792
rect 16807 10761 16819 10764
rect 16761 10755 16819 10761
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 17494 10752 17500 10804
rect 17552 10792 17558 10804
rect 21085 10795 21143 10801
rect 21085 10792 21097 10795
rect 17552 10764 21097 10792
rect 17552 10752 17558 10764
rect 21085 10761 21097 10764
rect 21131 10761 21143 10795
rect 22370 10792 22376 10804
rect 21085 10755 21143 10761
rect 22066 10764 22376 10792
rect 16666 10724 16672 10736
rect 11256 10696 16672 10724
rect 8573 10659 8631 10665
rect 8573 10656 8585 10659
rect 7892 10628 8585 10656
rect 7892 10616 7898 10628
rect 8573 10625 8585 10628
rect 8619 10625 8631 10659
rect 8573 10619 8631 10625
rect 11149 10659 11207 10665
rect 11149 10625 11161 10659
rect 11195 10625 11207 10659
rect 11149 10619 11207 10625
rect 1228 10588 1256 10616
rect 1765 10591 1823 10597
rect 1765 10588 1777 10591
rect 1228 10560 1777 10588
rect 1765 10557 1777 10560
rect 1811 10557 1823 10591
rect 1765 10551 1823 10557
rect 3160 10529 3188 10616
rect 4246 10548 4252 10600
rect 4304 10588 4310 10600
rect 4801 10591 4859 10597
rect 4801 10588 4813 10591
rect 4304 10560 4813 10588
rect 4304 10548 4310 10560
rect 4801 10557 4813 10560
rect 4847 10557 4859 10591
rect 11057 10591 11115 10597
rect 11057 10588 11069 10591
rect 4801 10551 4859 10557
rect 6196 10560 11069 10588
rect 6196 10529 6224 10560
rect 11057 10557 11069 10560
rect 11103 10557 11115 10591
rect 11057 10551 11115 10557
rect 3145 10523 3203 10529
rect 3145 10489 3157 10523
rect 3191 10489 3203 10523
rect 3145 10483 3203 10489
rect 6181 10523 6239 10529
rect 6181 10489 6193 10523
rect 6227 10489 6239 10523
rect 6181 10483 6239 10489
rect 6641 10523 6699 10529
rect 6641 10489 6653 10523
rect 6687 10520 6699 10523
rect 11256 10520 11284 10696
rect 16666 10684 16672 10696
rect 16724 10684 16730 10736
rect 17954 10724 17960 10736
rect 16868 10696 17960 10724
rect 11606 10616 11612 10668
rect 11664 10616 11670 10668
rect 13469 10659 13527 10665
rect 13469 10625 13481 10659
rect 13515 10656 13527 10659
rect 13630 10656 13636 10668
rect 13515 10628 13636 10656
rect 13515 10625 13527 10628
rect 13469 10619 13527 10625
rect 13630 10616 13636 10628
rect 13688 10616 13694 10668
rect 13722 10616 13728 10668
rect 13780 10616 13786 10668
rect 13814 10616 13820 10668
rect 13872 10656 13878 10668
rect 14366 10665 14372 10668
rect 14001 10659 14059 10665
rect 14001 10656 14013 10659
rect 13872 10628 14013 10656
rect 13872 10616 13878 10628
rect 14001 10625 14013 10628
rect 14047 10625 14059 10659
rect 14360 10656 14372 10665
rect 14327 10628 14372 10656
rect 14001 10619 14059 10625
rect 14360 10619 14372 10628
rect 14366 10616 14372 10619
rect 14424 10616 14430 10668
rect 14642 10616 14648 10668
rect 14700 10656 14706 10668
rect 15565 10659 15623 10665
rect 15565 10656 15577 10659
rect 14700 10628 15577 10656
rect 14700 10616 14706 10628
rect 15565 10625 15577 10628
rect 15611 10625 15623 10659
rect 15565 10619 15623 10625
rect 16114 10616 16120 10668
rect 16172 10656 16178 10668
rect 16868 10665 16896 10696
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 18414 10684 18420 10736
rect 18472 10724 18478 10736
rect 18966 10724 18972 10736
rect 18472 10696 18972 10724
rect 18472 10684 18478 10696
rect 18966 10684 18972 10696
rect 19024 10724 19030 10736
rect 19024 10696 21404 10724
rect 19024 10684 19030 10696
rect 21376 10668 21404 10696
rect 16301 10659 16359 10665
rect 16301 10656 16313 10659
rect 16172 10628 16313 10656
rect 16172 10616 16178 10628
rect 16301 10625 16313 10628
rect 16347 10625 16359 10659
rect 16301 10619 16359 10625
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 18785 10659 18843 10665
rect 18785 10625 18797 10659
rect 18831 10656 18843 10659
rect 19426 10656 19432 10668
rect 18831 10628 19432 10656
rect 18831 10625 18843 10628
rect 18785 10619 18843 10625
rect 12253 10591 12311 10597
rect 12253 10557 12265 10591
rect 12299 10557 12311 10591
rect 12253 10551 12311 10557
rect 6687 10492 11284 10520
rect 11333 10523 11391 10529
rect 6687 10489 6699 10492
rect 6641 10483 6699 10489
rect 11333 10489 11345 10523
rect 11379 10520 11391 10523
rect 11514 10520 11520 10532
rect 11379 10492 11520 10520
rect 11379 10489 11391 10492
rect 11333 10483 11391 10489
rect 11514 10480 11520 10492
rect 11572 10480 11578 10532
rect 12268 10520 12296 10551
rect 14090 10548 14096 10600
rect 14148 10548 14154 10600
rect 16574 10548 16580 10600
rect 16632 10588 16638 10600
rect 17052 10588 17080 10619
rect 19426 10616 19432 10628
rect 19484 10616 19490 10668
rect 20001 10659 20059 10665
rect 20001 10625 20013 10659
rect 20047 10656 20059 10659
rect 20047 10628 20392 10656
rect 20047 10625 20059 10628
rect 20001 10619 20059 10625
rect 16632 10560 17080 10588
rect 16632 10548 16638 10560
rect 17218 10548 17224 10600
rect 17276 10588 17282 10600
rect 20257 10591 20315 10597
rect 17276 10560 19196 10588
rect 17276 10548 17282 10560
rect 12345 10523 12403 10529
rect 12345 10520 12357 10523
rect 12268 10492 12357 10520
rect 12345 10489 12357 10492
rect 12391 10489 12403 10523
rect 12345 10483 12403 10489
rect 1673 10455 1731 10461
rect 1673 10421 1685 10455
rect 1719 10452 1731 10455
rect 5074 10452 5080 10464
rect 1719 10424 5080 10452
rect 1719 10421 1731 10424
rect 1673 10415 1731 10421
rect 5074 10412 5080 10424
rect 5132 10412 5138 10464
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 7009 10455 7067 10461
rect 7009 10452 7021 10455
rect 6972 10424 7021 10452
rect 6972 10412 6978 10424
rect 7009 10421 7021 10424
rect 7055 10421 7067 10455
rect 7009 10415 7067 10421
rect 10045 10455 10103 10461
rect 10045 10421 10057 10455
rect 10091 10452 10103 10455
rect 10318 10452 10324 10464
rect 10091 10424 10324 10452
rect 10091 10421 10103 10424
rect 10045 10415 10103 10421
rect 10318 10412 10324 10424
rect 10376 10412 10382 10464
rect 10410 10412 10416 10464
rect 10468 10412 10474 10464
rect 12526 10412 12532 10464
rect 12584 10452 12590 10464
rect 13909 10455 13967 10461
rect 13909 10452 13921 10455
rect 12584 10424 13921 10452
rect 12584 10412 12590 10424
rect 13909 10421 13921 10424
rect 13955 10421 13967 10455
rect 14108 10452 14136 10548
rect 16393 10523 16451 10529
rect 16393 10489 16405 10523
rect 16439 10520 16451 10523
rect 19058 10520 19064 10532
rect 16439 10492 19064 10520
rect 16439 10489 16451 10492
rect 16393 10483 16451 10489
rect 19058 10480 19064 10492
rect 19116 10480 19122 10532
rect 19168 10520 19196 10560
rect 20257 10557 20269 10591
rect 20303 10557 20315 10591
rect 20364 10588 20392 10628
rect 20438 10616 20444 10668
rect 20496 10656 20502 10668
rect 21269 10659 21327 10665
rect 21269 10656 21281 10659
rect 20496 10628 21281 10656
rect 20496 10616 20502 10628
rect 21269 10625 21281 10628
rect 21315 10625 21327 10659
rect 21269 10619 21327 10625
rect 21358 10616 21364 10668
rect 21416 10616 21422 10668
rect 21910 10616 21916 10668
rect 21968 10656 21974 10668
rect 22066 10656 22094 10764
rect 22370 10752 22376 10764
rect 22428 10752 22434 10804
rect 22922 10752 22928 10804
rect 22980 10752 22986 10804
rect 23014 10752 23020 10804
rect 23072 10792 23078 10804
rect 23385 10795 23443 10801
rect 23385 10792 23397 10795
rect 23072 10764 23397 10792
rect 23072 10752 23078 10764
rect 23385 10761 23397 10764
rect 23431 10761 23443 10795
rect 23385 10755 23443 10761
rect 22940 10665 22968 10752
rect 21968 10628 22094 10656
rect 22934 10659 22992 10665
rect 21968 10616 21974 10628
rect 22934 10625 22946 10659
rect 22980 10625 22992 10659
rect 22934 10619 22992 10625
rect 23198 10616 23204 10668
rect 23256 10616 23262 10668
rect 23293 10659 23351 10665
rect 23293 10625 23305 10659
rect 23339 10625 23351 10659
rect 23293 10619 23351 10625
rect 20898 10588 20904 10600
rect 20364 10560 20904 10588
rect 20257 10551 20315 10557
rect 20272 10520 20300 10551
rect 20898 10548 20904 10560
rect 20956 10548 20962 10600
rect 20993 10591 21051 10597
rect 20993 10557 21005 10591
rect 21039 10588 21051 10591
rect 21039 10560 21588 10588
rect 21039 10557 21051 10560
rect 20993 10551 21051 10557
rect 21453 10523 21511 10529
rect 21453 10520 21465 10523
rect 19168 10492 19334 10520
rect 20272 10492 21465 10520
rect 14458 10452 14464 10464
rect 14108 10424 14464 10452
rect 13909 10415 13967 10421
rect 14458 10412 14464 10424
rect 14516 10412 14522 10464
rect 18877 10455 18935 10461
rect 18877 10421 18889 10455
rect 18923 10452 18935 10455
rect 19150 10452 19156 10464
rect 18923 10424 19156 10452
rect 18923 10421 18935 10424
rect 18877 10415 18935 10421
rect 19150 10412 19156 10424
rect 19208 10412 19214 10464
rect 19306 10452 19334 10492
rect 21453 10489 21465 10492
rect 21499 10489 21511 10523
rect 21560 10520 21588 10560
rect 21634 10548 21640 10600
rect 21692 10588 21698 10600
rect 21692 10560 22094 10588
rect 21692 10548 21698 10560
rect 21821 10523 21879 10529
rect 21821 10520 21833 10523
rect 21560 10492 21833 10520
rect 21453 10483 21511 10489
rect 21821 10489 21833 10492
rect 21867 10489 21879 10523
rect 21821 10483 21879 10489
rect 20349 10455 20407 10461
rect 20349 10452 20361 10455
rect 19306 10424 20361 10452
rect 20349 10421 20361 10424
rect 20395 10421 20407 10455
rect 22066 10452 22094 10560
rect 23308 10452 23336 10619
rect 22066 10424 23336 10452
rect 20349 10415 20407 10421
rect 1104 10362 23828 10384
rect 1104 10310 1918 10362
rect 1970 10310 1982 10362
rect 2034 10310 2046 10362
rect 2098 10310 2110 10362
rect 2162 10310 2174 10362
rect 2226 10310 2238 10362
rect 2290 10310 7918 10362
rect 7970 10310 7982 10362
rect 8034 10310 8046 10362
rect 8098 10310 8110 10362
rect 8162 10310 8174 10362
rect 8226 10310 8238 10362
rect 8290 10310 13918 10362
rect 13970 10310 13982 10362
rect 14034 10310 14046 10362
rect 14098 10310 14110 10362
rect 14162 10310 14174 10362
rect 14226 10310 14238 10362
rect 14290 10310 19918 10362
rect 19970 10310 19982 10362
rect 20034 10310 20046 10362
rect 20098 10310 20110 10362
rect 20162 10310 20174 10362
rect 20226 10310 20238 10362
rect 20290 10310 23828 10362
rect 1104 10288 23828 10310
rect 1578 10208 1584 10260
rect 1636 10248 1642 10260
rect 2498 10248 2504 10260
rect 1636 10220 2504 10248
rect 1636 10208 1642 10220
rect 2498 10208 2504 10220
rect 2556 10248 2562 10260
rect 5997 10251 6055 10257
rect 2556 10220 4016 10248
rect 2556 10208 2562 10220
rect 3510 10180 3516 10192
rect 1596 10152 3516 10180
rect 1596 10121 1624 10152
rect 3510 10140 3516 10152
rect 3568 10140 3574 10192
rect 3605 10183 3663 10189
rect 3605 10149 3617 10183
rect 3651 10180 3663 10183
rect 3878 10180 3884 10192
rect 3651 10152 3884 10180
rect 3651 10149 3663 10152
rect 3605 10143 3663 10149
rect 3878 10140 3884 10152
rect 3936 10140 3942 10192
rect 3988 10121 4016 10220
rect 5997 10217 6009 10251
rect 6043 10248 6055 10251
rect 6362 10248 6368 10260
rect 6043 10220 6368 10248
rect 6043 10217 6055 10220
rect 5997 10211 6055 10217
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 8113 10251 8171 10257
rect 8113 10248 8125 10251
rect 7248 10220 8125 10248
rect 7248 10208 7254 10220
rect 8113 10217 8125 10220
rect 8159 10217 8171 10251
rect 8113 10211 8171 10217
rect 12253 10251 12311 10257
rect 12253 10217 12265 10251
rect 12299 10248 12311 10251
rect 12299 10220 13492 10248
rect 12299 10217 12311 10220
rect 12253 10211 12311 10217
rect 7742 10140 7748 10192
rect 7800 10180 7806 10192
rect 9125 10183 9183 10189
rect 7800 10152 7972 10180
rect 7800 10140 7806 10152
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10081 1639 10115
rect 3973 10115 4031 10121
rect 1581 10075 1639 10081
rect 2746 10084 3004 10112
rect 2222 10004 2228 10056
rect 2280 10044 2286 10056
rect 2590 10044 2596 10056
rect 2280 10016 2596 10044
rect 2280 10004 2286 10016
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 2133 9979 2191 9985
rect 2133 9945 2145 9979
rect 2179 9976 2191 9979
rect 2746 9976 2774 10084
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10013 2927 10047
rect 2869 10007 2927 10013
rect 2179 9948 2774 9976
rect 2179 9945 2191 9948
rect 2133 9939 2191 9945
rect 1302 9868 1308 9920
rect 1360 9908 1366 9920
rect 2225 9911 2283 9917
rect 2225 9908 2237 9911
rect 1360 9880 2237 9908
rect 1360 9868 1366 9880
rect 2225 9877 2237 9880
rect 2271 9877 2283 9911
rect 2884 9908 2912 10007
rect 2976 9976 3004 10084
rect 3973 10081 3985 10115
rect 4019 10081 4031 10115
rect 3973 10075 4031 10081
rect 4338 10072 4344 10124
rect 4396 10072 4402 10124
rect 7834 10112 7840 10124
rect 5736 10084 7840 10112
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10044 3111 10047
rect 4356 10044 4384 10072
rect 5736 10053 5764 10084
rect 7834 10072 7840 10084
rect 7892 10072 7898 10124
rect 3099 10016 4384 10044
rect 5721 10047 5779 10053
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 5721 10013 5733 10047
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 7944 10044 7972 10152
rect 9125 10149 9137 10183
rect 9171 10180 9183 10183
rect 10594 10180 10600 10192
rect 9171 10152 10600 10180
rect 9171 10149 9183 10152
rect 9125 10143 9183 10149
rect 10594 10140 10600 10152
rect 10652 10140 10658 10192
rect 13464 10180 13492 10220
rect 13630 10208 13636 10260
rect 13688 10248 13694 10260
rect 13909 10251 13967 10257
rect 13909 10248 13921 10251
rect 13688 10220 13921 10248
rect 13688 10208 13694 10220
rect 13909 10217 13921 10220
rect 13955 10217 13967 10251
rect 13909 10211 13967 10217
rect 15657 10251 15715 10257
rect 15657 10217 15669 10251
rect 15703 10248 15715 10251
rect 17770 10248 17776 10260
rect 15703 10220 17776 10248
rect 15703 10217 15715 10220
rect 15657 10211 15715 10217
rect 17770 10208 17776 10220
rect 17828 10208 17834 10260
rect 20346 10248 20352 10260
rect 18524 10220 20352 10248
rect 13464 10152 14228 10180
rect 14200 10124 14228 10152
rect 8757 10115 8815 10121
rect 8757 10081 8769 10115
rect 8803 10112 8815 10115
rect 9858 10112 9864 10124
rect 8803 10084 9864 10112
rect 8803 10081 8815 10084
rect 8757 10075 8815 10081
rect 9858 10072 9864 10084
rect 9916 10072 9922 10124
rect 11146 10072 11152 10124
rect 11204 10112 11210 10124
rect 11204 10084 12112 10112
rect 11204 10072 11210 10084
rect 11532 10056 11560 10084
rect 9493 10047 9551 10053
rect 9493 10044 9505 10047
rect 7944 10016 9505 10044
rect 4522 9976 4528 9988
rect 2976 9948 4528 9976
rect 4522 9936 4528 9948
rect 4580 9936 4586 9988
rect 5534 9976 5540 9988
rect 4632 9948 5540 9976
rect 4632 9908 4660 9948
rect 5534 9936 5540 9948
rect 5592 9936 5598 9988
rect 5920 9976 5948 10007
rect 5994 9976 6000 9988
rect 5920 9948 6000 9976
rect 5994 9936 6000 9948
rect 6052 9936 6058 9988
rect 7944 9985 7972 10016
rect 9493 10013 9505 10016
rect 9539 10013 9551 10047
rect 9493 10007 9551 10013
rect 6181 9979 6239 9985
rect 6181 9945 6193 9979
rect 6227 9945 6239 9979
rect 6181 9939 6239 9945
rect 7929 9979 7987 9985
rect 7929 9945 7941 9979
rect 7975 9945 7987 9979
rect 7929 9939 7987 9945
rect 2884 9880 4660 9908
rect 2225 9871 2283 9877
rect 4706 9868 4712 9920
rect 4764 9908 4770 9920
rect 6196 9908 6224 9939
rect 9306 9936 9312 9988
rect 9364 9976 9370 9988
rect 9401 9979 9459 9985
rect 9401 9976 9413 9979
rect 9364 9948 9413 9976
rect 9364 9936 9370 9948
rect 9401 9945 9413 9948
rect 9447 9945 9459 9979
rect 9508 9976 9536 10007
rect 11514 10004 11520 10056
rect 11572 10004 11578 10056
rect 11790 10004 11796 10056
rect 11848 10044 11854 10056
rect 12084 10053 12112 10084
rect 14182 10072 14188 10124
rect 14240 10072 14246 10124
rect 18524 10121 18552 10220
rect 20346 10208 20352 10220
rect 20404 10208 20410 10260
rect 20625 10251 20683 10257
rect 20625 10217 20637 10251
rect 20671 10248 20683 10251
rect 20671 10220 21772 10248
rect 20671 10217 20683 10220
rect 20625 10211 20683 10217
rect 18785 10183 18843 10189
rect 18785 10149 18797 10183
rect 18831 10180 18843 10183
rect 18874 10180 18880 10192
rect 18831 10152 18880 10180
rect 18831 10149 18843 10152
rect 18785 10143 18843 10149
rect 18874 10140 18880 10152
rect 18932 10140 18938 10192
rect 18509 10115 18567 10121
rect 18509 10081 18521 10115
rect 18555 10081 18567 10115
rect 18509 10075 18567 10081
rect 11885 10047 11943 10053
rect 11885 10044 11897 10047
rect 11848 10016 11897 10044
rect 11848 10004 11854 10016
rect 11885 10013 11897 10016
rect 11931 10013 11943 10047
rect 11885 10007 11943 10013
rect 12069 10047 12127 10053
rect 12069 10013 12081 10047
rect 12115 10013 12127 10047
rect 12069 10007 12127 10013
rect 12526 10004 12532 10056
rect 12584 10004 12590 10056
rect 12802 10053 12808 10056
rect 12796 10007 12808 10053
rect 12860 10044 12866 10056
rect 12860 10016 12896 10044
rect 12802 10004 12808 10007
rect 12860 10004 12866 10016
rect 15562 10004 15568 10056
rect 15620 10004 15626 10056
rect 17037 10047 17095 10053
rect 17037 10013 17049 10047
rect 17083 10044 17095 10047
rect 19245 10047 19303 10053
rect 19245 10044 19257 10047
rect 17083 10016 19257 10044
rect 17083 10013 17095 10016
rect 17037 10007 17095 10013
rect 19245 10013 19257 10016
rect 19291 10044 19303 10047
rect 19334 10044 19340 10056
rect 19291 10016 19340 10044
rect 19291 10013 19303 10016
rect 19245 10007 19303 10013
rect 19334 10004 19340 10016
rect 19392 10044 19398 10056
rect 20070 10044 20076 10056
rect 19392 10016 20076 10044
rect 19392 10004 19398 10016
rect 20070 10004 20076 10016
rect 20128 10004 20134 10056
rect 20717 10047 20775 10053
rect 20717 10013 20729 10047
rect 20763 10044 20775 10047
rect 21450 10044 21456 10056
rect 20763 10016 21456 10044
rect 20763 10013 20775 10016
rect 20717 10007 20775 10013
rect 21450 10004 21456 10016
rect 21508 10004 21514 10056
rect 21744 10044 21772 10220
rect 23290 10072 23296 10124
rect 23348 10072 23354 10124
rect 22002 10044 22008 10056
rect 21744 10016 22008 10044
rect 22002 10004 22008 10016
rect 22060 10004 22066 10056
rect 22189 10047 22247 10053
rect 22189 10044 22201 10047
rect 22112 10016 22201 10044
rect 12618 9976 12624 9988
rect 9508 9948 12624 9976
rect 9401 9939 9459 9945
rect 12618 9936 12624 9948
rect 12676 9936 12682 9988
rect 14090 9936 14096 9988
rect 14148 9976 14154 9988
rect 15298 9979 15356 9985
rect 15298 9976 15310 9979
rect 14148 9948 15310 9976
rect 14148 9936 14154 9948
rect 15298 9945 15310 9948
rect 15344 9945 15356 9979
rect 15298 9939 15356 9945
rect 16792 9979 16850 9985
rect 16792 9945 16804 9979
rect 16838 9976 16850 9979
rect 17586 9976 17592 9988
rect 16838 9948 17592 9976
rect 16838 9945 16850 9948
rect 16792 9939 16850 9945
rect 17586 9936 17592 9948
rect 17644 9936 17650 9988
rect 18138 9936 18144 9988
rect 18196 9936 18202 9988
rect 18230 9936 18236 9988
rect 18288 9985 18294 9988
rect 18288 9939 18300 9985
rect 18288 9936 18294 9939
rect 18506 9936 18512 9988
rect 18564 9976 18570 9988
rect 19061 9979 19119 9985
rect 19061 9976 19073 9979
rect 18564 9948 19073 9976
rect 18564 9936 18570 9948
rect 19061 9945 19073 9948
rect 19107 9945 19119 9979
rect 19061 9939 19119 9945
rect 19150 9936 19156 9988
rect 19208 9976 19214 9988
rect 19490 9979 19548 9985
rect 19490 9976 19502 9979
rect 19208 9948 19502 9976
rect 19208 9936 19214 9948
rect 19490 9945 19502 9948
rect 19536 9945 19548 9979
rect 19490 9939 19548 9945
rect 20984 9979 21042 9985
rect 20984 9945 20996 9979
rect 21030 9976 21042 9979
rect 21910 9976 21916 9988
rect 21030 9948 21916 9976
rect 21030 9945 21042 9948
rect 20984 9939 21042 9945
rect 21910 9936 21916 9948
rect 21968 9936 21974 9988
rect 6270 9908 6276 9920
rect 4764 9880 6276 9908
rect 4764 9868 4770 9880
rect 6270 9868 6276 9880
rect 6328 9868 6334 9920
rect 8478 9868 8484 9920
rect 8536 9908 8542 9920
rect 8941 9911 8999 9917
rect 8941 9908 8953 9911
rect 8536 9880 8953 9908
rect 8536 9868 8542 9880
rect 8941 9877 8953 9880
rect 8987 9877 8999 9911
rect 8941 9871 8999 9877
rect 10686 9868 10692 9920
rect 10744 9908 10750 9920
rect 10781 9911 10839 9917
rect 10781 9908 10793 9911
rect 10744 9880 10793 9908
rect 10744 9868 10750 9880
rect 10781 9877 10793 9880
rect 10827 9877 10839 9911
rect 10781 9871 10839 9877
rect 11333 9911 11391 9917
rect 11333 9877 11345 9911
rect 11379 9908 11391 9911
rect 11606 9908 11612 9920
rect 11379 9880 11612 9908
rect 11379 9877 11391 9880
rect 11333 9871 11391 9877
rect 11606 9868 11612 9880
rect 11664 9868 11670 9920
rect 12526 9868 12532 9920
rect 12584 9908 12590 9920
rect 14185 9911 14243 9917
rect 14185 9908 14197 9911
rect 12584 9880 14197 9908
rect 12584 9868 12590 9880
rect 14185 9877 14197 9880
rect 14231 9877 14243 9911
rect 14185 9871 14243 9877
rect 17126 9868 17132 9920
rect 17184 9868 17190 9920
rect 18156 9908 18184 9936
rect 18601 9911 18659 9917
rect 18601 9908 18613 9911
rect 18156 9880 18613 9908
rect 18601 9877 18613 9880
rect 18647 9877 18659 9911
rect 18601 9871 18659 9877
rect 20898 9868 20904 9920
rect 20956 9908 20962 9920
rect 21634 9908 21640 9920
rect 20956 9880 21640 9908
rect 20956 9868 20962 9880
rect 21634 9868 21640 9880
rect 21692 9868 21698 9920
rect 22112 9917 22140 10016
rect 22189 10013 22201 10016
rect 22235 10013 22247 10047
rect 22189 10007 22247 10013
rect 22462 10004 22468 10056
rect 22520 10004 22526 10056
rect 22738 10004 22744 10056
rect 22796 10044 22802 10056
rect 22833 10047 22891 10053
rect 22833 10044 22845 10047
rect 22796 10016 22845 10044
rect 22796 10004 22802 10016
rect 22833 10013 22845 10016
rect 22879 10013 22891 10047
rect 22833 10007 22891 10013
rect 22097 9911 22155 9917
rect 22097 9877 22109 9911
rect 22143 9877 22155 9911
rect 22097 9871 22155 9877
rect 1104 9818 23828 9840
rect 1104 9766 2658 9818
rect 2710 9766 2722 9818
rect 2774 9766 2786 9818
rect 2838 9766 2850 9818
rect 2902 9766 2914 9818
rect 2966 9766 2978 9818
rect 3030 9766 8658 9818
rect 8710 9766 8722 9818
rect 8774 9766 8786 9818
rect 8838 9766 8850 9818
rect 8902 9766 8914 9818
rect 8966 9766 8978 9818
rect 9030 9766 14658 9818
rect 14710 9766 14722 9818
rect 14774 9766 14786 9818
rect 14838 9766 14850 9818
rect 14902 9766 14914 9818
rect 14966 9766 14978 9818
rect 15030 9766 20658 9818
rect 20710 9766 20722 9818
rect 20774 9766 20786 9818
rect 20838 9766 20850 9818
rect 20902 9766 20914 9818
rect 20966 9766 20978 9818
rect 21030 9766 23828 9818
rect 1104 9744 23828 9766
rect 2222 9704 2228 9716
rect 2148 9676 2228 9704
rect 2148 9645 2176 9676
rect 2222 9664 2228 9676
rect 2280 9664 2286 9716
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 6730 9704 6736 9716
rect 6052 9676 6736 9704
rect 6052 9664 6058 9676
rect 6730 9664 6736 9676
rect 6788 9704 6794 9716
rect 10318 9704 10324 9716
rect 6788 9676 10324 9704
rect 6788 9664 6794 9676
rect 10318 9664 10324 9676
rect 10376 9704 10382 9716
rect 14366 9704 14372 9716
rect 10376 9676 14372 9704
rect 10376 9664 10382 9676
rect 14366 9664 14372 9676
rect 14424 9664 14430 9716
rect 14458 9664 14464 9716
rect 14516 9704 14522 9716
rect 14516 9676 14688 9704
rect 14516 9664 14522 9676
rect 14660 9648 14688 9676
rect 21358 9664 21364 9716
rect 21416 9704 21422 9716
rect 21416 9676 21680 9704
rect 21416 9664 21422 9676
rect 21652 9674 21680 9676
rect 2133 9639 2191 9645
rect 2133 9605 2145 9639
rect 2179 9605 2191 9639
rect 2133 9599 2191 9605
rect 3326 9596 3332 9648
rect 3384 9636 3390 9648
rect 6365 9639 6423 9645
rect 6365 9636 6377 9639
rect 3384 9608 6377 9636
rect 3384 9596 3390 9608
rect 6365 9605 6377 9608
rect 6411 9605 6423 9639
rect 6365 9599 6423 9605
rect 6822 9596 6828 9648
rect 6880 9636 6886 9648
rect 11974 9636 11980 9648
rect 6880 9608 11980 9636
rect 6880 9596 6886 9608
rect 11974 9596 11980 9608
rect 12032 9596 12038 9648
rect 13940 9639 13998 9645
rect 13940 9605 13952 9639
rect 13986 9636 13998 9639
rect 14274 9636 14280 9648
rect 13986 9608 14280 9636
rect 13986 9605 13998 9608
rect 13940 9599 13998 9605
rect 14274 9596 14280 9608
rect 14332 9596 14338 9648
rect 14642 9596 14648 9648
rect 14700 9596 14706 9648
rect 15470 9596 15476 9648
rect 15528 9636 15534 9648
rect 16390 9636 16396 9648
rect 15528 9608 16396 9636
rect 15528 9596 15534 9608
rect 16390 9596 16396 9608
rect 16448 9596 16454 9648
rect 16666 9596 16672 9648
rect 16724 9596 16730 9648
rect 19518 9596 19524 9648
rect 19576 9636 19582 9648
rect 21652 9646 21772 9674
rect 19622 9639 19680 9645
rect 19622 9636 19634 9639
rect 19576 9608 19634 9636
rect 19576 9596 19582 9608
rect 19622 9605 19634 9608
rect 19668 9605 19680 9639
rect 21094 9639 21152 9645
rect 21094 9636 21106 9639
rect 19622 9599 19680 9605
rect 20824 9608 21106 9636
rect 20824 9580 20852 9608
rect 21094 9605 21106 9608
rect 21140 9605 21152 9639
rect 21744 9636 21772 9646
rect 21744 9608 21864 9636
rect 21094 9599 21152 9605
rect 2222 9528 2228 9580
rect 2280 9528 2286 9580
rect 2685 9571 2743 9577
rect 2685 9537 2697 9571
rect 2731 9568 2743 9571
rect 3237 9571 3295 9577
rect 2731 9540 3188 9568
rect 2731 9537 2743 9540
rect 2685 9531 2743 9537
rect 1581 9503 1639 9509
rect 1581 9469 1593 9503
rect 1627 9500 1639 9503
rect 2958 9500 2964 9512
rect 1627 9472 2964 9500
rect 1627 9469 1639 9472
rect 1581 9463 1639 9469
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 3160 9500 3188 9540
rect 3237 9537 3249 9571
rect 3283 9568 3295 9571
rect 4154 9568 4160 9580
rect 3283 9540 4160 9568
rect 3283 9537 3295 9540
rect 3237 9531 3295 9537
rect 4154 9528 4160 9540
rect 4212 9528 4218 9580
rect 4453 9571 4511 9577
rect 4453 9537 4465 9571
rect 4499 9568 4511 9571
rect 4614 9568 4620 9580
rect 4499 9540 4620 9568
rect 4499 9537 4511 9540
rect 4453 9531 4511 9537
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 4706 9528 4712 9580
rect 4764 9528 4770 9580
rect 5074 9577 5080 9580
rect 5057 9571 5080 9577
rect 5057 9537 5069 9571
rect 5057 9531 5080 9537
rect 5074 9528 5080 9531
rect 5132 9528 5138 9580
rect 5534 9528 5540 9580
rect 5592 9568 5598 9580
rect 8113 9571 8171 9577
rect 5592 9540 5856 9568
rect 5592 9528 5598 9540
rect 3602 9500 3608 9512
rect 3160 9472 3608 9500
rect 3602 9460 3608 9472
rect 3660 9460 3666 9512
rect 4798 9460 4804 9512
rect 4856 9460 4862 9512
rect 5828 9500 5856 9540
rect 8113 9537 8125 9571
rect 8159 9568 8171 9571
rect 10410 9568 10416 9580
rect 8159 9540 8340 9568
rect 8159 9537 8171 9540
rect 8113 9531 8171 9537
rect 8205 9503 8263 9509
rect 8205 9500 8217 9503
rect 5828 9472 8217 9500
rect 8205 9469 8217 9472
rect 8251 9469 8263 9503
rect 8205 9463 8263 9469
rect 2406 9392 2412 9444
rect 2464 9392 2470 9444
rect 2590 9392 2596 9444
rect 2648 9432 2654 9444
rect 7098 9432 7104 9444
rect 2648 9404 3464 9432
rect 2648 9392 2654 9404
rect 3234 9324 3240 9376
rect 3292 9364 3298 9376
rect 3329 9367 3387 9373
rect 3329 9364 3341 9367
rect 3292 9336 3341 9364
rect 3292 9324 3298 9336
rect 3329 9333 3341 9336
rect 3375 9333 3387 9367
rect 3436 9364 3464 9404
rect 5736 9404 7104 9432
rect 5736 9364 5764 9404
rect 7098 9392 7104 9404
rect 7156 9392 7162 9444
rect 3436 9336 5764 9364
rect 6181 9367 6239 9373
rect 3329 9327 3387 9333
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 7190 9364 7196 9376
rect 6227 9336 7196 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 8312 9364 8340 9540
rect 8404 9540 10416 9568
rect 8404 9441 8432 9540
rect 10410 9528 10416 9540
rect 10468 9528 10474 9580
rect 10505 9571 10563 9577
rect 10505 9537 10517 9571
rect 10551 9537 10563 9571
rect 10505 9531 10563 9537
rect 8665 9503 8723 9509
rect 8665 9469 8677 9503
rect 8711 9500 8723 9503
rect 9306 9500 9312 9512
rect 8711 9472 9312 9500
rect 8711 9469 8723 9472
rect 8665 9463 8723 9469
rect 9306 9460 9312 9472
rect 9364 9460 9370 9512
rect 8389 9435 8447 9441
rect 8389 9401 8401 9435
rect 8435 9401 8447 9435
rect 9324 9432 9352 9460
rect 10520 9432 10548 9531
rect 10594 9528 10600 9580
rect 10652 9528 10658 9580
rect 11514 9528 11520 9580
rect 11572 9568 11578 9580
rect 11793 9571 11851 9577
rect 11793 9568 11805 9571
rect 11572 9540 11805 9568
rect 11572 9528 11578 9540
rect 11793 9537 11805 9540
rect 11839 9537 11851 9571
rect 11793 9531 11851 9537
rect 13446 9528 13452 9580
rect 13504 9568 13510 9580
rect 14090 9568 14096 9580
rect 13504 9540 14096 9568
rect 13504 9528 13510 9540
rect 14090 9528 14096 9540
rect 14148 9528 14154 9580
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9568 14519 9571
rect 19889 9571 19947 9577
rect 14507 9540 17448 9568
rect 14507 9537 14519 9540
rect 14461 9531 14519 9537
rect 11241 9503 11299 9509
rect 11241 9469 11253 9503
rect 11287 9500 11299 9503
rect 11698 9500 11704 9512
rect 11287 9472 11704 9500
rect 11287 9469 11299 9472
rect 11241 9463 11299 9469
rect 11698 9460 11704 9472
rect 11756 9460 11762 9512
rect 12526 9460 12532 9512
rect 12584 9460 12590 9512
rect 14185 9503 14243 9509
rect 14185 9469 14197 9503
rect 14231 9500 14243 9503
rect 14369 9503 14427 9509
rect 14369 9500 14381 9503
rect 14231 9472 14381 9500
rect 14231 9469 14243 9472
rect 14185 9463 14243 9469
rect 14369 9469 14381 9472
rect 14415 9469 14427 9503
rect 14369 9463 14427 9469
rect 12986 9432 12992 9444
rect 9324 9404 9444 9432
rect 10520 9404 12992 9432
rect 8389 9395 8447 9401
rect 9217 9367 9275 9373
rect 9217 9364 9229 9367
rect 8312 9336 9229 9364
rect 9217 9333 9229 9336
rect 9263 9364 9275 9367
rect 9306 9364 9312 9376
rect 9263 9336 9312 9364
rect 9263 9333 9275 9336
rect 9217 9327 9275 9333
rect 9306 9324 9312 9336
rect 9364 9324 9370 9376
rect 9416 9364 9444 9404
rect 12986 9392 12992 9404
rect 13044 9392 13050 9444
rect 17420 9376 17448 9540
rect 19889 9537 19901 9571
rect 19935 9537 19947 9571
rect 19889 9531 19947 9537
rect 17862 9392 17868 9444
rect 17920 9432 17926 9444
rect 18509 9435 18567 9441
rect 18509 9432 18521 9435
rect 17920 9404 18521 9432
rect 17920 9392 17926 9404
rect 18509 9401 18521 9404
rect 18555 9401 18567 9435
rect 18509 9395 18567 9401
rect 9674 9364 9680 9376
rect 9416 9336 9680 9364
rect 9674 9324 9680 9336
rect 9732 9364 9738 9376
rect 11238 9364 11244 9376
rect 9732 9336 11244 9364
rect 9732 9324 9738 9336
rect 11238 9324 11244 9336
rect 11296 9364 11302 9376
rect 11609 9367 11667 9373
rect 11609 9364 11621 9367
rect 11296 9336 11621 9364
rect 11296 9324 11302 9336
rect 11609 9333 11621 9336
rect 11655 9333 11667 9367
rect 11609 9327 11667 9333
rect 11882 9324 11888 9376
rect 11940 9364 11946 9376
rect 11977 9367 12035 9373
rect 11977 9364 11989 9367
rect 11940 9336 11989 9364
rect 11940 9324 11946 9336
rect 11977 9333 11989 9336
rect 12023 9333 12035 9367
rect 11977 9327 12035 9333
rect 12802 9324 12808 9376
rect 12860 9324 12866 9376
rect 14182 9324 14188 9376
rect 14240 9364 14246 9376
rect 15378 9364 15384 9376
rect 14240 9336 15384 9364
rect 14240 9324 14246 9336
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 17402 9324 17408 9376
rect 17460 9324 17466 9376
rect 17954 9324 17960 9376
rect 18012 9324 18018 9376
rect 19904 9364 19932 9531
rect 20806 9528 20812 9580
rect 20864 9528 20870 9580
rect 21453 9572 21511 9577
rect 21836 9574 21864 9608
rect 21652 9572 21864 9574
rect 21453 9571 21864 9572
rect 21453 9537 21465 9571
rect 21499 9546 21864 9571
rect 21499 9544 21680 9546
rect 21499 9537 21511 9544
rect 21453 9531 21511 9537
rect 21910 9528 21916 9580
rect 21968 9568 21974 9580
rect 22077 9571 22135 9577
rect 22077 9568 22089 9571
rect 21968 9540 22089 9568
rect 21968 9528 21974 9540
rect 22077 9537 22089 9540
rect 22123 9537 22135 9571
rect 22077 9531 22135 9537
rect 23474 9528 23480 9580
rect 23532 9528 23538 9580
rect 21358 9509 21364 9512
rect 21354 9500 21364 9509
rect 21319 9472 21364 9500
rect 21354 9463 21364 9472
rect 21358 9460 21364 9463
rect 21416 9460 21422 9512
rect 21726 9460 21732 9512
rect 21784 9500 21790 9512
rect 21821 9503 21879 9509
rect 21821 9500 21833 9503
rect 21784 9472 21833 9500
rect 21784 9460 21790 9472
rect 21821 9469 21833 9472
rect 21867 9469 21879 9503
rect 21821 9463 21879 9469
rect 19981 9435 20039 9441
rect 19981 9401 19993 9435
rect 20027 9432 20039 9435
rect 20346 9432 20352 9444
rect 20027 9404 20352 9432
rect 20027 9401 20039 9404
rect 19981 9395 20039 9401
rect 20346 9392 20352 9404
rect 20404 9392 20410 9444
rect 21545 9435 21603 9441
rect 21545 9401 21557 9435
rect 21591 9401 21603 9435
rect 21545 9395 21603 9401
rect 21560 9364 21588 9395
rect 23290 9392 23296 9444
rect 23348 9392 23354 9444
rect 19904 9336 21588 9364
rect 23106 9324 23112 9376
rect 23164 9364 23170 9376
rect 23201 9367 23259 9373
rect 23201 9364 23213 9367
rect 23164 9336 23213 9364
rect 23164 9324 23170 9336
rect 23201 9333 23213 9336
rect 23247 9333 23259 9367
rect 23201 9327 23259 9333
rect 1104 9274 23828 9296
rect 1104 9222 1918 9274
rect 1970 9222 1982 9274
rect 2034 9222 2046 9274
rect 2098 9222 2110 9274
rect 2162 9222 2174 9274
rect 2226 9222 2238 9274
rect 2290 9222 7918 9274
rect 7970 9222 7982 9274
rect 8034 9222 8046 9274
rect 8098 9222 8110 9274
rect 8162 9222 8174 9274
rect 8226 9222 8238 9274
rect 8290 9222 13918 9274
rect 13970 9222 13982 9274
rect 14034 9222 14046 9274
rect 14098 9222 14110 9274
rect 14162 9222 14174 9274
rect 14226 9222 14238 9274
rect 14290 9222 19918 9274
rect 19970 9222 19982 9274
rect 20034 9222 20046 9274
rect 20098 9222 20110 9274
rect 20162 9222 20174 9274
rect 20226 9222 20238 9274
rect 20290 9222 23828 9274
rect 1104 9200 23828 9222
rect 2133 9163 2191 9169
rect 2133 9129 2145 9163
rect 2179 9160 2191 9163
rect 5074 9160 5080 9172
rect 2179 9132 5080 9160
rect 2179 9129 2191 9132
rect 2133 9123 2191 9129
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 8386 9120 8392 9172
rect 8444 9160 8450 9172
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 8444 9132 9045 9160
rect 8444 9120 8450 9132
rect 9033 9129 9045 9132
rect 9079 9129 9091 9163
rect 9033 9123 9091 9129
rect 9858 9120 9864 9172
rect 9916 9160 9922 9172
rect 10597 9163 10655 9169
rect 10597 9160 10609 9163
rect 9916 9132 10609 9160
rect 9916 9120 9922 9132
rect 10597 9129 10609 9132
rect 10643 9129 10655 9163
rect 10597 9123 10655 9129
rect 11974 9120 11980 9172
rect 12032 9120 12038 9172
rect 12526 9120 12532 9172
rect 12584 9120 12590 9172
rect 12802 9120 12808 9172
rect 12860 9160 12866 9172
rect 12860 9132 17356 9160
rect 12860 9120 12866 9132
rect 9214 9092 9220 9104
rect 8772 9064 9220 9092
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8956 1639 8959
rect 2130 8956 2136 8968
rect 1627 8928 2136 8956
rect 1627 8925 1639 8928
rect 1581 8919 1639 8925
rect 2130 8916 2136 8928
rect 2188 8916 2194 8968
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 2271 8928 2774 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 1854 8848 1860 8900
rect 1912 8888 1918 8900
rect 2470 8891 2528 8897
rect 2470 8888 2482 8891
rect 1912 8860 2482 8888
rect 1912 8848 1918 8860
rect 2470 8857 2482 8860
rect 2516 8857 2528 8891
rect 2746 8888 2774 8928
rect 2958 8916 2964 8968
rect 3016 8956 3022 8968
rect 3510 8956 3516 8968
rect 3016 8928 3516 8956
rect 3016 8916 3022 8928
rect 3510 8916 3516 8928
rect 3568 8916 3574 8968
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8956 3847 8959
rect 3970 8956 3976 8968
rect 3835 8928 3976 8956
rect 3835 8925 3847 8928
rect 3789 8919 3847 8925
rect 3970 8916 3976 8928
rect 4028 8916 4034 8968
rect 4062 8916 4068 8968
rect 4120 8916 4126 8968
rect 4706 8956 4712 8968
rect 4172 8928 4712 8956
rect 4172 8888 4200 8928
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 5074 8916 5080 8968
rect 5132 8956 5138 8968
rect 8478 8956 8484 8968
rect 5132 8928 8484 8956
rect 5132 8916 5138 8928
rect 8478 8916 8484 8928
rect 8536 8916 8542 8968
rect 8772 8965 8800 9064
rect 9214 9052 9220 9064
rect 9272 9052 9278 9104
rect 17328 9092 17356 9132
rect 17402 9120 17408 9172
rect 17460 9160 17466 9172
rect 19150 9160 19156 9172
rect 17460 9132 19156 9160
rect 17460 9120 17466 9132
rect 19150 9120 19156 9132
rect 19208 9160 19214 9172
rect 19208 9132 23336 9160
rect 19208 9120 19214 9132
rect 18417 9095 18475 9101
rect 17328 9064 18368 9092
rect 17586 8984 17592 9036
rect 17644 9024 17650 9036
rect 17773 9027 17831 9033
rect 17773 9024 17785 9027
rect 17644 8996 17785 9024
rect 17644 8984 17650 8996
rect 17773 8993 17785 8996
rect 17819 8993 17831 9027
rect 18340 9024 18368 9064
rect 18417 9061 18429 9095
rect 18463 9092 18475 9095
rect 18598 9092 18604 9104
rect 18463 9064 18604 9092
rect 18463 9061 18475 9064
rect 18417 9055 18475 9061
rect 18598 9052 18604 9064
rect 18656 9052 18662 9104
rect 18877 9095 18935 9101
rect 18877 9061 18889 9095
rect 18923 9092 18935 9095
rect 19242 9092 19248 9104
rect 18923 9064 19248 9092
rect 18923 9061 18935 9064
rect 18877 9055 18935 9061
rect 19242 9052 19248 9064
rect 19300 9052 19306 9104
rect 20346 9052 20352 9104
rect 20404 9052 20410 9104
rect 20530 9052 20536 9104
rect 20588 9092 20594 9104
rect 20625 9095 20683 9101
rect 20625 9092 20637 9095
rect 20588 9064 20637 9092
rect 20588 9052 20594 9064
rect 20625 9061 20637 9064
rect 20671 9061 20683 9095
rect 20625 9055 20683 9061
rect 18340 8996 19380 9024
rect 17773 8987 17831 8993
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8925 8815 8959
rect 8757 8919 8815 8925
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 4338 8897 4344 8900
rect 2746 8860 4200 8888
rect 2470 8851 2528 8857
rect 4332 8851 4344 8897
rect 4338 8848 4344 8851
rect 4396 8848 4402 8900
rect 5626 8888 5632 8900
rect 5072 8860 5632 8888
rect 3602 8780 3608 8832
rect 3660 8780 3666 8832
rect 3973 8823 4031 8829
rect 3973 8789 3985 8823
rect 4019 8820 4031 8823
rect 5072 8820 5100 8860
rect 5626 8848 5632 8860
rect 5684 8848 5690 8900
rect 7009 8891 7067 8897
rect 7009 8857 7021 8891
rect 7055 8857 7067 8891
rect 7009 8851 7067 8857
rect 4019 8792 5100 8820
rect 4019 8789 4031 8792
rect 3973 8783 4031 8789
rect 5442 8780 5448 8832
rect 5500 8780 5506 8832
rect 6546 8780 6552 8832
rect 6604 8820 6610 8832
rect 7024 8820 7052 8851
rect 8570 8848 8576 8900
rect 8628 8888 8634 8900
rect 9140 8888 9168 8919
rect 9214 8916 9220 8968
rect 9272 8916 9278 8968
rect 9306 8916 9312 8968
rect 9364 8956 9370 8968
rect 10689 8959 10747 8965
rect 10689 8956 10701 8959
rect 9364 8928 10701 8956
rect 9364 8916 9370 8928
rect 10689 8925 10701 8928
rect 10735 8925 10747 8959
rect 10689 8919 10747 8925
rect 13814 8916 13820 8968
rect 13872 8916 13878 8968
rect 13906 8916 13912 8968
rect 13964 8916 13970 8968
rect 14182 8916 14188 8968
rect 14240 8956 14246 8968
rect 15841 8959 15899 8965
rect 14240 8928 14688 8956
rect 14240 8916 14246 8928
rect 8628 8860 9168 8888
rect 8628 8848 8634 8860
rect 6604 8792 7052 8820
rect 9140 8820 9168 8860
rect 9484 8891 9542 8897
rect 9484 8857 9496 8891
rect 9530 8888 9542 8891
rect 9858 8888 9864 8900
rect 9530 8860 9864 8888
rect 9530 8857 9542 8860
rect 9484 8851 9542 8857
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 13538 8848 13544 8900
rect 13596 8888 13602 8900
rect 13642 8891 13700 8897
rect 13642 8888 13654 8891
rect 13596 8860 13654 8888
rect 13596 8848 13602 8860
rect 13642 8857 13654 8860
rect 13688 8857 13700 8891
rect 13832 8888 13860 8916
rect 14093 8891 14151 8897
rect 14093 8888 14105 8891
rect 13832 8860 14105 8888
rect 13642 8851 13700 8857
rect 14093 8857 14105 8860
rect 14139 8888 14151 8891
rect 14550 8888 14556 8900
rect 14139 8860 14556 8888
rect 14139 8857 14151 8860
rect 14093 8851 14151 8857
rect 14550 8848 14556 8860
rect 14608 8848 14614 8900
rect 14660 8888 14688 8928
rect 15841 8925 15853 8959
rect 15887 8956 15899 8959
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 15887 8928 18000 8956
rect 15887 8925 15899 8928
rect 15841 8919 15899 8925
rect 17972 8900 18000 8928
rect 18064 8928 19257 8956
rect 15933 8891 15991 8897
rect 15933 8888 15945 8891
rect 14660 8860 15945 8888
rect 15933 8857 15945 8860
rect 15979 8857 15991 8891
rect 15933 8851 15991 8857
rect 17954 8848 17960 8900
rect 18012 8848 18018 8900
rect 10226 8820 10232 8832
rect 9140 8792 10232 8820
rect 6604 8780 6610 8792
rect 10226 8780 10232 8792
rect 10284 8780 10290 8832
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 14642 8820 14648 8832
rect 13872 8792 14648 8820
rect 13872 8780 13878 8792
rect 14642 8780 14648 8792
rect 14700 8820 14706 8832
rect 18064 8820 18092 8928
rect 19245 8925 19257 8928
rect 19291 8925 19303 8959
rect 19352 8956 19380 8996
rect 19352 8928 19656 8956
rect 19245 8919 19303 8925
rect 18506 8848 18512 8900
rect 18564 8848 18570 8900
rect 18690 8848 18696 8900
rect 18748 8888 18754 8900
rect 19490 8891 19548 8897
rect 19490 8888 19502 8891
rect 18748 8860 19502 8888
rect 18748 8848 18754 8860
rect 19490 8857 19502 8860
rect 19536 8857 19548 8891
rect 19490 8851 19548 8857
rect 14700 8792 18092 8820
rect 14700 8780 14706 8792
rect 18782 8780 18788 8832
rect 18840 8820 18846 8832
rect 18969 8823 19027 8829
rect 18969 8820 18981 8823
rect 18840 8792 18981 8820
rect 18840 8780 18846 8792
rect 18969 8789 18981 8792
rect 19015 8789 19027 8823
rect 19628 8820 19656 8928
rect 20364 8888 20392 9052
rect 22646 8984 22652 9036
rect 22704 9024 22710 9036
rect 23109 9027 23167 9033
rect 23109 9024 23121 9027
rect 22704 8996 23121 9024
rect 22704 8984 22710 8996
rect 23109 8993 23121 8996
rect 23155 8993 23167 9027
rect 23109 8987 23167 8993
rect 20717 8959 20775 8965
rect 20717 8925 20729 8959
rect 20763 8956 20775 8959
rect 21358 8956 21364 8968
rect 20763 8928 21364 8956
rect 20763 8925 20775 8928
rect 20717 8919 20775 8925
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 22833 8959 22891 8965
rect 22833 8956 22845 8959
rect 22066 8928 22845 8956
rect 20962 8891 21020 8897
rect 20962 8888 20974 8891
rect 20364 8860 20974 8888
rect 20962 8857 20974 8860
rect 21008 8857 21020 8891
rect 22066 8888 22094 8928
rect 22833 8925 22845 8928
rect 22879 8925 22891 8959
rect 22833 8919 22891 8925
rect 20962 8851 21020 8857
rect 21100 8860 22094 8888
rect 21100 8820 21128 8860
rect 23308 8832 23336 9132
rect 19628 8792 21128 8820
rect 18969 8783 19027 8789
rect 22094 8780 22100 8832
rect 22152 8780 22158 8832
rect 23290 8780 23296 8832
rect 23348 8780 23354 8832
rect 1104 8730 23828 8752
rect 1104 8678 2658 8730
rect 2710 8678 2722 8730
rect 2774 8678 2786 8730
rect 2838 8678 2850 8730
rect 2902 8678 2914 8730
rect 2966 8678 2978 8730
rect 3030 8678 8658 8730
rect 8710 8678 8722 8730
rect 8774 8678 8786 8730
rect 8838 8678 8850 8730
rect 8902 8678 8914 8730
rect 8966 8678 8978 8730
rect 9030 8678 14658 8730
rect 14710 8678 14722 8730
rect 14774 8678 14786 8730
rect 14838 8678 14850 8730
rect 14902 8678 14914 8730
rect 14966 8678 14978 8730
rect 15030 8678 20658 8730
rect 20710 8678 20722 8730
rect 20774 8678 20786 8730
rect 20838 8678 20850 8730
rect 20902 8678 20914 8730
rect 20966 8678 20978 8730
rect 21030 8678 23828 8730
rect 1104 8656 23828 8678
rect 1673 8619 1731 8625
rect 1673 8585 1685 8619
rect 1719 8616 1731 8619
rect 9214 8616 9220 8628
rect 1719 8588 9220 8616
rect 1719 8585 1731 8588
rect 1673 8579 1731 8585
rect 9214 8576 9220 8588
rect 9272 8576 9278 8628
rect 13906 8576 13912 8628
rect 13964 8616 13970 8628
rect 14369 8619 14427 8625
rect 14369 8616 14381 8619
rect 13964 8588 14381 8616
rect 13964 8576 13970 8588
rect 14369 8585 14381 8588
rect 14415 8585 14427 8619
rect 15286 8616 15292 8628
rect 14369 8579 14427 8585
rect 14568 8588 15292 8616
rect 2498 8548 2504 8560
rect 1780 8520 2504 8548
rect 1780 8489 1808 8520
rect 2498 8508 2504 8520
rect 2556 8548 2562 8560
rect 3326 8548 3332 8560
rect 2556 8520 3332 8548
rect 2556 8508 2562 8520
rect 3326 8508 3332 8520
rect 3384 8508 3390 8560
rect 3602 8557 3608 8560
rect 3596 8548 3608 8557
rect 3563 8520 3608 8548
rect 3596 8511 3608 8520
rect 3602 8508 3608 8511
rect 3660 8508 3666 8560
rect 3694 8508 3700 8560
rect 3752 8508 3758 8560
rect 3970 8508 3976 8560
rect 4028 8508 4034 8560
rect 5166 8508 5172 8560
rect 5224 8548 5230 8560
rect 6365 8551 6423 8557
rect 6365 8548 6377 8551
rect 5224 8520 6377 8548
rect 5224 8508 5230 8520
rect 6365 8517 6377 8520
rect 6411 8517 6423 8551
rect 6365 8511 6423 8517
rect 7190 8508 7196 8560
rect 7248 8508 7254 8560
rect 7834 8508 7840 8560
rect 7892 8548 7898 8560
rect 7929 8551 7987 8557
rect 7929 8548 7941 8551
rect 7892 8520 7941 8548
rect 7892 8508 7898 8520
rect 7929 8517 7941 8520
rect 7975 8517 7987 8551
rect 7929 8511 7987 8517
rect 9401 8551 9459 8557
rect 9401 8517 9413 8551
rect 9447 8548 9459 8551
rect 9674 8548 9680 8560
rect 9447 8520 9680 8548
rect 9447 8517 9459 8520
rect 9401 8511 9459 8517
rect 9674 8508 9680 8520
rect 9732 8508 9738 8560
rect 11333 8551 11391 8557
rect 11333 8517 11345 8551
rect 11379 8548 11391 8551
rect 14182 8548 14188 8560
rect 11379 8520 14188 8548
rect 11379 8517 11391 8520
rect 11333 8511 11391 8517
rect 14182 8508 14188 8520
rect 14240 8508 14246 8560
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8449 1823 8483
rect 1765 8443 1823 8449
rect 1854 8440 1860 8492
rect 1912 8440 1918 8492
rect 2130 8440 2136 8492
rect 2188 8440 2194 8492
rect 2981 8483 3039 8489
rect 2981 8449 2993 8483
rect 3027 8480 3039 8483
rect 3712 8480 3740 8508
rect 3027 8452 3740 8480
rect 3988 8480 4016 8508
rect 5534 8480 5540 8492
rect 3988 8452 5540 8480
rect 3027 8449 3039 8452
rect 2981 8443 3039 8449
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 5925 8483 5983 8489
rect 5925 8449 5937 8483
rect 5971 8480 5983 8483
rect 7208 8480 7236 8508
rect 8205 8483 8263 8489
rect 8205 8480 8217 8483
rect 5971 8452 7144 8480
rect 7208 8452 8217 8480
rect 5971 8449 5983 8452
rect 5925 8443 5983 8449
rect 1872 8353 1900 8440
rect 1857 8347 1915 8353
rect 1857 8313 1869 8347
rect 1903 8313 1915 8347
rect 2148 8344 2176 8440
rect 3234 8372 3240 8424
rect 3292 8372 3298 8424
rect 3326 8372 3332 8424
rect 3384 8372 3390 8424
rect 4356 8384 4844 8412
rect 4356 8344 4384 8384
rect 2148 8316 2360 8344
rect 1857 8307 1915 8313
rect 2332 8276 2360 8316
rect 4264 8316 4384 8344
rect 4816 8344 4844 8384
rect 6178 8372 6184 8424
rect 6236 8372 6242 8424
rect 7116 8412 7144 8452
rect 8205 8449 8217 8452
rect 8251 8449 8263 8483
rect 8205 8443 8263 8449
rect 12434 8440 12440 8492
rect 12492 8440 12498 8492
rect 14461 8486 14519 8489
rect 14568 8486 14596 8588
rect 15286 8576 15292 8588
rect 15344 8616 15350 8628
rect 16114 8616 16120 8628
rect 15344 8588 16120 8616
rect 15344 8576 15350 8588
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 16206 8576 16212 8628
rect 16264 8576 16270 8628
rect 19058 8576 19064 8628
rect 19116 8616 19122 8628
rect 19245 8619 19303 8625
rect 19245 8616 19257 8619
rect 19116 8588 19257 8616
rect 19116 8576 19122 8588
rect 19245 8585 19257 8588
rect 19291 8616 19303 8619
rect 21266 8616 21272 8628
rect 19291 8588 21272 8616
rect 19291 8585 19303 8588
rect 19245 8579 19303 8585
rect 21266 8576 21272 8588
rect 21324 8576 21330 8628
rect 21361 8619 21419 8625
rect 21361 8585 21373 8619
rect 21407 8616 21419 8619
rect 21818 8616 21824 8628
rect 21407 8588 21824 8616
rect 21407 8585 21419 8588
rect 21361 8579 21419 8585
rect 21818 8576 21824 8588
rect 21876 8576 21882 8628
rect 22186 8576 22192 8628
rect 22244 8616 22250 8628
rect 23201 8619 23259 8625
rect 23201 8616 23213 8619
rect 22244 8588 23213 8616
rect 22244 8576 22250 8588
rect 23201 8585 23213 8588
rect 23247 8585 23259 8619
rect 23201 8579 23259 8585
rect 17405 8551 17463 8557
rect 17405 8548 17417 8551
rect 15396 8520 17417 8548
rect 15396 8492 15424 8520
rect 17405 8517 17417 8520
rect 17451 8548 17463 8551
rect 18506 8548 18512 8560
rect 17451 8520 18512 8548
rect 17451 8517 17463 8520
rect 17405 8511 17463 8517
rect 18506 8508 18512 8520
rect 18564 8508 18570 8560
rect 20530 8508 20536 8560
rect 20588 8548 20594 8560
rect 20910 8551 20968 8557
rect 20910 8548 20922 8551
rect 20588 8520 20922 8548
rect 20588 8508 20594 8520
rect 20910 8517 20922 8520
rect 20956 8517 20968 8551
rect 23385 8551 23443 8557
rect 23385 8548 23397 8551
rect 20910 8511 20968 8517
rect 21192 8520 23397 8548
rect 14461 8483 14596 8486
rect 14461 8449 14473 8483
rect 14507 8458 14596 8483
rect 14507 8449 14519 8458
rect 14461 8443 14519 8449
rect 15378 8440 15384 8492
rect 15436 8440 15442 8492
rect 15746 8440 15752 8492
rect 15804 8489 15810 8492
rect 15804 8443 15816 8489
rect 15804 8440 15810 8443
rect 16298 8440 16304 8492
rect 16356 8440 16362 8492
rect 16761 8483 16819 8489
rect 16761 8449 16773 8483
rect 16807 8480 16819 8483
rect 17126 8480 17132 8492
rect 16807 8452 17132 8480
rect 16807 8449 16819 8452
rect 16761 8443 16819 8449
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 17313 8483 17371 8489
rect 17313 8449 17325 8483
rect 17359 8480 17371 8483
rect 17359 8452 17908 8480
rect 17359 8449 17371 8452
rect 17313 8443 17371 8449
rect 8938 8412 8944 8424
rect 7116 8384 8944 8412
rect 8938 8372 8944 8384
rect 8996 8372 9002 8424
rect 11793 8415 11851 8421
rect 11793 8381 11805 8415
rect 11839 8412 11851 8415
rect 13722 8412 13728 8424
rect 11839 8384 13728 8412
rect 11839 8381 11851 8384
rect 11793 8375 11851 8381
rect 13722 8372 13728 8384
rect 13780 8372 13786 8424
rect 15010 8412 15016 8424
rect 14476 8384 15016 8412
rect 8849 8347 8907 8353
rect 4816 8316 5304 8344
rect 3510 8276 3516 8288
rect 2332 8248 3516 8276
rect 3510 8236 3516 8248
rect 3568 8236 3574 8288
rect 3602 8236 3608 8288
rect 3660 8276 3666 8288
rect 4264 8276 4292 8316
rect 3660 8248 4292 8276
rect 3660 8236 3666 8248
rect 4522 8236 4528 8288
rect 4580 8276 4586 8288
rect 4709 8279 4767 8285
rect 4709 8276 4721 8279
rect 4580 8248 4721 8276
rect 4580 8236 4586 8248
rect 4709 8245 4721 8248
rect 4755 8245 4767 8279
rect 4709 8239 4767 8245
rect 4801 8279 4859 8285
rect 4801 8245 4813 8279
rect 4847 8276 4859 8279
rect 4890 8276 4896 8288
rect 4847 8248 4896 8276
rect 4847 8245 4859 8248
rect 4801 8239 4859 8245
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 5276 8276 5304 8316
rect 8849 8313 8861 8347
rect 8895 8344 8907 8347
rect 9033 8347 9091 8353
rect 9033 8344 9045 8347
rect 8895 8316 9045 8344
rect 8895 8313 8907 8316
rect 8849 8307 8907 8313
rect 9033 8313 9045 8316
rect 9079 8313 9091 8347
rect 9033 8307 9091 8313
rect 12345 8347 12403 8353
rect 12345 8313 12357 8347
rect 12391 8344 12403 8347
rect 14476 8344 14504 8384
rect 15010 8372 15016 8384
rect 15068 8372 15074 8424
rect 16025 8415 16083 8421
rect 16025 8381 16037 8415
rect 16071 8412 16083 8415
rect 16574 8412 16580 8424
rect 16071 8384 16580 8412
rect 16071 8381 16083 8384
rect 16025 8375 16083 8381
rect 16574 8372 16580 8384
rect 16632 8372 16638 8424
rect 17880 8412 17908 8452
rect 17954 8440 17960 8492
rect 18012 8440 18018 8492
rect 20438 8480 20444 8492
rect 20180 8452 20444 8480
rect 18874 8412 18880 8424
rect 17880 8384 18880 8412
rect 18874 8372 18880 8384
rect 18932 8372 18938 8424
rect 19794 8372 19800 8424
rect 19852 8372 19858 8424
rect 12391 8316 14504 8344
rect 14645 8347 14703 8353
rect 12391 8313 12403 8316
rect 12345 8307 12403 8313
rect 14645 8313 14657 8347
rect 14691 8344 14703 8347
rect 14691 8316 15148 8344
rect 14691 8313 14703 8316
rect 14645 8307 14703 8313
rect 5902 8276 5908 8288
rect 5276 8248 5908 8276
rect 5902 8236 5908 8248
rect 5960 8236 5966 8288
rect 6454 8236 6460 8288
rect 6512 8276 6518 8288
rect 8941 8279 8999 8285
rect 8941 8276 8953 8279
rect 6512 8248 8953 8276
rect 6512 8236 6518 8248
rect 8941 8245 8953 8248
rect 8987 8245 8999 8279
rect 8941 8239 8999 8245
rect 10042 8236 10048 8288
rect 10100 8236 10106 8288
rect 15120 8276 15148 8316
rect 16114 8304 16120 8356
rect 16172 8344 16178 8356
rect 16666 8344 16672 8356
rect 16172 8316 16672 8344
rect 16172 8304 16178 8316
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 17773 8347 17831 8353
rect 17773 8313 17785 8347
rect 17819 8313 17831 8347
rect 17773 8307 17831 8313
rect 17865 8347 17923 8353
rect 17865 8313 17877 8347
rect 17911 8344 17923 8347
rect 18230 8344 18236 8356
rect 17911 8316 18236 8344
rect 17911 8313 17923 8316
rect 17865 8307 17923 8313
rect 16390 8276 16396 8288
rect 15120 8248 16396 8276
rect 16390 8236 16396 8248
rect 16448 8236 16454 8288
rect 17788 8276 17816 8307
rect 18230 8304 18236 8316
rect 18288 8304 18294 8356
rect 19812 8344 19840 8372
rect 20180 8344 20208 8452
rect 20438 8440 20444 8452
rect 20496 8480 20502 8492
rect 21192 8489 21220 8520
rect 23385 8517 23397 8520
rect 23431 8517 23443 8551
rect 23385 8511 23443 8517
rect 21177 8483 21235 8489
rect 20496 8452 21128 8480
rect 20496 8440 20502 8452
rect 21100 8412 21128 8452
rect 21177 8449 21189 8483
rect 21223 8449 21235 8483
rect 21177 8443 21235 8449
rect 21269 8483 21327 8489
rect 21269 8449 21281 8483
rect 21315 8480 21327 8483
rect 21634 8480 21640 8492
rect 21315 8452 21640 8480
rect 21315 8449 21327 8452
rect 21269 8443 21327 8449
rect 21634 8440 21640 8452
rect 21692 8440 21698 8492
rect 21726 8440 21732 8492
rect 21784 8480 21790 8492
rect 21821 8483 21879 8489
rect 21821 8480 21833 8483
rect 21784 8452 21833 8480
rect 21784 8440 21790 8452
rect 21821 8449 21833 8452
rect 21867 8449 21879 8483
rect 22077 8483 22135 8489
rect 22077 8480 22089 8483
rect 21821 8443 21879 8449
rect 21928 8452 22089 8480
rect 21928 8412 21956 8452
rect 22077 8449 22089 8452
rect 22123 8449 22135 8483
rect 22077 8443 22135 8449
rect 23290 8440 23296 8492
rect 23348 8440 23354 8492
rect 21100 8384 21956 8412
rect 18340 8316 19840 8344
rect 19904 8316 20208 8344
rect 18340 8276 18368 8316
rect 17788 8248 18368 8276
rect 19797 8279 19855 8285
rect 19797 8245 19809 8279
rect 19843 8276 19855 8279
rect 19904 8276 19932 8316
rect 19843 8248 19932 8276
rect 19843 8245 19855 8248
rect 19797 8239 19855 8245
rect 21174 8236 21180 8288
rect 21232 8276 21238 8288
rect 22462 8276 22468 8288
rect 21232 8248 22468 8276
rect 21232 8236 21238 8248
rect 22462 8236 22468 8248
rect 22520 8236 22526 8288
rect 1104 8186 23828 8208
rect 1104 8134 1918 8186
rect 1970 8134 1982 8186
rect 2034 8134 2046 8186
rect 2098 8134 2110 8186
rect 2162 8134 2174 8186
rect 2226 8134 2238 8186
rect 2290 8134 7918 8186
rect 7970 8134 7982 8186
rect 8034 8134 8046 8186
rect 8098 8134 8110 8186
rect 8162 8134 8174 8186
rect 8226 8134 8238 8186
rect 8290 8134 13918 8186
rect 13970 8134 13982 8186
rect 14034 8134 14046 8186
rect 14098 8134 14110 8186
rect 14162 8134 14174 8186
rect 14226 8134 14238 8186
rect 14290 8134 19918 8186
rect 19970 8134 19982 8186
rect 20034 8134 20046 8186
rect 20098 8134 20110 8186
rect 20162 8134 20174 8186
rect 20226 8134 20238 8186
rect 20290 8134 23828 8186
rect 1104 8112 23828 8134
rect 2222 8032 2228 8084
rect 2280 8072 2286 8084
rect 2406 8072 2412 8084
rect 2280 8044 2412 8072
rect 2280 8032 2286 8044
rect 2406 8032 2412 8044
rect 2464 8032 2470 8084
rect 3510 8032 3516 8084
rect 3568 8032 3574 8084
rect 3602 8032 3608 8084
rect 3660 8032 3666 8084
rect 3973 8075 4031 8081
rect 3973 8041 3985 8075
rect 4019 8072 4031 8075
rect 5166 8072 5172 8084
rect 4019 8044 5172 8072
rect 4019 8041 4031 8044
rect 3973 8035 4031 8041
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 8938 8032 8944 8084
rect 8996 8032 9002 8084
rect 9398 8032 9404 8084
rect 9456 8072 9462 8084
rect 12253 8075 12311 8081
rect 12253 8072 12265 8075
rect 9456 8044 12265 8072
rect 9456 8032 9462 8044
rect 12253 8041 12265 8044
rect 12299 8041 12311 8075
rect 12253 8035 12311 8041
rect 14274 8032 14280 8084
rect 14332 8072 14338 8084
rect 14458 8072 14464 8084
rect 14332 8044 14464 8072
rect 14332 8032 14338 8044
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 16390 8032 16396 8084
rect 16448 8072 16454 8084
rect 16448 8044 19840 8072
rect 16448 8032 16454 8044
rect 3528 8004 3556 8032
rect 4065 8007 4123 8013
rect 4065 8004 4077 8007
rect 3528 7976 4077 8004
rect 4065 7973 4077 7976
rect 4111 7973 4123 8007
rect 4065 7967 4123 7973
rect 10413 8007 10471 8013
rect 10413 7973 10425 8007
rect 10459 8004 10471 8007
rect 10502 8004 10508 8016
rect 10459 7976 10508 8004
rect 10459 7973 10471 7976
rect 10413 7967 10471 7973
rect 10502 7964 10508 7976
rect 10560 7964 10566 8016
rect 11974 7964 11980 8016
rect 12032 8004 12038 8016
rect 12032 7976 12434 8004
rect 12032 7964 12038 7976
rect 10686 7936 10692 7948
rect 3712 7908 3924 7936
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7837 1639 7871
rect 1581 7831 1639 7837
rect 2225 7871 2283 7877
rect 2225 7837 2237 7871
rect 2271 7868 2283 7871
rect 2314 7868 2320 7880
rect 2271 7840 2320 7868
rect 2271 7837 2283 7840
rect 2225 7831 2283 7837
rect 1596 7800 1624 7831
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 3712 7868 3740 7908
rect 2424 7840 3740 7868
rect 2424 7800 2452 7840
rect 3786 7828 3792 7880
rect 3844 7828 3850 7880
rect 3896 7868 3924 7908
rect 10336 7908 10692 7936
rect 4890 7868 4896 7880
rect 3896 7840 4896 7868
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 5442 7828 5448 7880
rect 5500 7828 5506 7880
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 1596 7772 2452 7800
rect 2492 7803 2550 7809
rect 2492 7769 2504 7803
rect 2538 7800 2550 7803
rect 2590 7800 2596 7812
rect 2538 7772 2596 7800
rect 2538 7769 2550 7772
rect 2492 7763 2550 7769
rect 2590 7760 2596 7772
rect 2648 7760 2654 7812
rect 3142 7760 3148 7812
rect 3200 7800 3206 7812
rect 4338 7800 4344 7812
rect 3200 7772 4344 7800
rect 3200 7760 3206 7772
rect 4338 7760 4344 7772
rect 4396 7760 4402 7812
rect 4982 7760 4988 7812
rect 5040 7800 5046 7812
rect 5178 7803 5236 7809
rect 5178 7800 5190 7803
rect 5040 7772 5190 7800
rect 5040 7760 5046 7772
rect 5178 7769 5190 7772
rect 5224 7769 5236 7803
rect 5178 7763 5236 7769
rect 5350 7760 5356 7812
rect 5408 7800 5414 7812
rect 5552 7800 5580 7831
rect 5626 7828 5632 7880
rect 5684 7868 5690 7880
rect 5793 7871 5851 7877
rect 5793 7868 5805 7871
rect 5684 7840 5805 7868
rect 5684 7828 5690 7840
rect 5793 7837 5805 7840
rect 5839 7837 5851 7871
rect 5793 7831 5851 7837
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7868 7435 7871
rect 7466 7868 7472 7880
rect 7423 7840 7472 7868
rect 7423 7837 7435 7840
rect 7377 7831 7435 7837
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 9490 7828 9496 7880
rect 9548 7868 9554 7880
rect 10336 7877 10364 7908
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 9548 7840 10333 7868
rect 9548 7828 9554 7840
rect 10321 7837 10333 7840
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 10597 7871 10655 7877
rect 10597 7837 10609 7871
rect 10643 7868 10655 7871
rect 10778 7868 10784 7880
rect 10643 7840 10784 7868
rect 10643 7837 10655 7840
rect 10597 7831 10655 7837
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 12158 7828 12164 7880
rect 12216 7828 12222 7880
rect 12406 7868 12434 7976
rect 19812 7945 19840 8044
rect 21358 8032 21364 8084
rect 21416 8072 21422 8084
rect 23201 8075 23259 8081
rect 23201 8072 23213 8075
rect 21416 8044 23213 8072
rect 21416 8032 21422 8044
rect 23201 8041 23213 8044
rect 23247 8041 23259 8075
rect 23201 8035 23259 8041
rect 19797 7939 19855 7945
rect 19797 7905 19809 7939
rect 19843 7905 19855 7939
rect 21818 7936 21824 7948
rect 19797 7899 19855 7905
rect 21468 7908 21824 7936
rect 13909 7871 13967 7877
rect 12406 7840 13768 7868
rect 7622 7803 7680 7809
rect 7622 7800 7634 7803
rect 5408 7772 5580 7800
rect 5644 7772 7634 7800
rect 5408 7760 5414 7772
rect 2133 7735 2191 7741
rect 2133 7701 2145 7735
rect 2179 7732 2191 7735
rect 5644 7732 5672 7772
rect 7622 7769 7634 7772
rect 7668 7769 7680 7803
rect 7622 7763 7680 7769
rect 9950 7760 9956 7812
rect 10008 7800 10014 7812
rect 10054 7803 10112 7809
rect 10054 7800 10066 7803
rect 10008 7772 10066 7800
rect 10008 7760 10014 7772
rect 10054 7769 10066 7772
rect 10100 7769 10112 7803
rect 10054 7763 10112 7769
rect 10956 7803 11014 7809
rect 10956 7769 10968 7803
rect 11002 7800 11014 7803
rect 12710 7800 12716 7812
rect 11002 7772 12716 7800
rect 11002 7769 11014 7772
rect 10956 7763 11014 7769
rect 12710 7760 12716 7772
rect 12768 7760 12774 7812
rect 13630 7760 13636 7812
rect 13688 7809 13694 7812
rect 13688 7763 13700 7809
rect 13740 7800 13768 7840
rect 13909 7837 13921 7871
rect 13955 7868 13967 7871
rect 14185 7871 14243 7877
rect 14185 7868 14197 7871
rect 13955 7840 14197 7868
rect 13955 7837 13967 7840
rect 13909 7831 13967 7837
rect 14185 7837 14197 7840
rect 14231 7837 14243 7871
rect 14185 7831 14243 7837
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7868 14335 7871
rect 14323 7840 14504 7868
rect 14323 7837 14335 7840
rect 14277 7831 14335 7837
rect 14476 7800 14504 7840
rect 15930 7828 15936 7880
rect 15988 7828 15994 7880
rect 16022 7828 16028 7880
rect 16080 7828 16086 7880
rect 16224 7840 18736 7868
rect 13740 7772 14504 7800
rect 13688 7760 13694 7763
rect 14476 7744 14504 7772
rect 15688 7803 15746 7809
rect 15688 7769 15700 7803
rect 15734 7800 15746 7803
rect 16224 7800 16252 7840
rect 16298 7809 16304 7812
rect 15734 7772 16252 7800
rect 15734 7769 15746 7772
rect 15688 7763 15746 7769
rect 16292 7763 16304 7809
rect 16298 7760 16304 7763
rect 16356 7760 16362 7812
rect 17678 7800 17684 7812
rect 17420 7772 17684 7800
rect 2179 7704 5672 7732
rect 6917 7735 6975 7741
rect 2179 7701 2191 7704
rect 2133 7695 2191 7701
rect 6917 7701 6929 7735
rect 6963 7732 6975 7735
rect 7834 7732 7840 7744
rect 6963 7704 7840 7732
rect 6963 7701 6975 7704
rect 6917 7695 6975 7701
rect 7834 7692 7840 7704
rect 7892 7692 7898 7744
rect 8757 7735 8815 7741
rect 8757 7701 8769 7735
rect 8803 7732 8815 7735
rect 10318 7732 10324 7744
rect 8803 7704 10324 7732
rect 8803 7701 8815 7704
rect 8757 7695 8815 7701
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 12066 7692 12072 7744
rect 12124 7692 12130 7744
rect 12529 7735 12587 7741
rect 12529 7701 12541 7735
rect 12575 7732 12587 7735
rect 14182 7732 14188 7744
rect 12575 7704 14188 7732
rect 12575 7701 12587 7704
rect 12529 7695 12587 7701
rect 14182 7692 14188 7704
rect 14240 7692 14246 7744
rect 14458 7692 14464 7744
rect 14516 7692 14522 7744
rect 14553 7735 14611 7741
rect 14553 7701 14565 7735
rect 14599 7732 14611 7735
rect 16114 7732 16120 7744
rect 14599 7704 16120 7732
rect 14599 7701 14611 7704
rect 14553 7695 14611 7701
rect 16114 7692 16120 7704
rect 16172 7692 16178 7744
rect 17420 7741 17448 7772
rect 17678 7760 17684 7772
rect 17736 7760 17742 7812
rect 18506 7760 18512 7812
rect 18564 7800 18570 7812
rect 18610 7803 18668 7809
rect 18610 7800 18622 7803
rect 18564 7772 18622 7800
rect 18564 7760 18570 7772
rect 18610 7769 18622 7772
rect 18656 7769 18668 7803
rect 18708 7800 18736 7840
rect 18874 7828 18880 7880
rect 18932 7828 18938 7880
rect 21468 7868 21496 7908
rect 21818 7896 21824 7908
rect 21876 7896 21882 7948
rect 22940 7908 23336 7936
rect 20180 7840 21496 7868
rect 19245 7803 19303 7809
rect 19245 7800 19257 7803
rect 18708 7772 19257 7800
rect 18610 7763 18668 7769
rect 19245 7769 19257 7772
rect 19291 7769 19303 7803
rect 19245 7763 19303 7769
rect 17405 7735 17463 7741
rect 17405 7701 17417 7735
rect 17451 7701 17463 7735
rect 17405 7695 17463 7701
rect 17497 7735 17555 7741
rect 17497 7701 17509 7735
rect 17543 7732 17555 7735
rect 18690 7732 18696 7744
rect 17543 7704 18696 7732
rect 17543 7701 17555 7704
rect 17497 7695 17555 7701
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 20180 7741 20208 7840
rect 21542 7828 21548 7880
rect 21600 7828 21606 7880
rect 21634 7828 21640 7880
rect 21692 7868 21698 7880
rect 22940 7868 22968 7908
rect 23308 7880 23336 7908
rect 21692 7840 22968 7868
rect 21692 7828 21698 7840
rect 23014 7828 23020 7880
rect 23072 7828 23078 7880
rect 23290 7828 23296 7880
rect 23348 7828 23354 7880
rect 21300 7803 21358 7809
rect 21300 7769 21312 7803
rect 21346 7800 21358 7803
rect 21726 7800 21732 7812
rect 21346 7772 21732 7800
rect 21346 7769 21358 7772
rect 21300 7763 21358 7769
rect 21726 7760 21732 7772
rect 21784 7760 21790 7812
rect 22738 7760 22744 7812
rect 22796 7809 22802 7812
rect 22796 7763 22808 7809
rect 22796 7760 22802 7763
rect 20165 7735 20223 7741
rect 20165 7701 20177 7735
rect 20211 7701 20223 7735
rect 20165 7695 20223 7701
rect 21174 7692 21180 7744
rect 21232 7732 21238 7744
rect 21637 7735 21695 7741
rect 21637 7732 21649 7735
rect 21232 7704 21649 7732
rect 21232 7692 21238 7704
rect 21637 7701 21649 7704
rect 21683 7701 21695 7735
rect 21637 7695 21695 7701
rect 1104 7642 23828 7664
rect 1104 7590 2658 7642
rect 2710 7590 2722 7642
rect 2774 7590 2786 7642
rect 2838 7590 2850 7642
rect 2902 7590 2914 7642
rect 2966 7590 2978 7642
rect 3030 7590 8658 7642
rect 8710 7590 8722 7642
rect 8774 7590 8786 7642
rect 8838 7590 8850 7642
rect 8902 7590 8914 7642
rect 8966 7590 8978 7642
rect 9030 7590 14658 7642
rect 14710 7590 14722 7642
rect 14774 7590 14786 7642
rect 14838 7590 14850 7642
rect 14902 7590 14914 7642
rect 14966 7590 14978 7642
rect 15030 7590 20658 7642
rect 20710 7590 20722 7642
rect 20774 7590 20786 7642
rect 20838 7590 20850 7642
rect 20902 7590 20914 7642
rect 20966 7590 20978 7642
rect 21030 7590 23828 7642
rect 1104 7568 23828 7590
rect 1670 7488 1676 7540
rect 1728 7488 1734 7540
rect 2222 7528 2228 7540
rect 1964 7500 2228 7528
rect 1688 7392 1716 7488
rect 1964 7404 1992 7500
rect 2222 7488 2228 7500
rect 2280 7488 2286 7540
rect 2409 7531 2467 7537
rect 2409 7497 2421 7531
rect 2455 7528 2467 7531
rect 3786 7528 3792 7540
rect 2455 7500 3792 7528
rect 2455 7497 2467 7500
rect 2409 7491 2467 7497
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 6086 7528 6092 7540
rect 4816 7500 6092 7528
rect 2041 7463 2099 7469
rect 2041 7429 2053 7463
rect 2087 7460 2099 7463
rect 3050 7460 3056 7472
rect 2087 7432 3056 7460
rect 2087 7429 2099 7432
rect 2041 7423 2099 7429
rect 3050 7420 3056 7432
rect 3108 7420 3114 7472
rect 3142 7420 3148 7472
rect 3200 7460 3206 7472
rect 3602 7469 3608 7472
rect 3237 7463 3295 7469
rect 3237 7460 3249 7463
rect 3200 7432 3249 7460
rect 3200 7420 3206 7432
rect 3237 7429 3249 7432
rect 3283 7429 3295 7463
rect 3237 7423 3295 7429
rect 3574 7463 3608 7469
rect 3574 7429 3586 7463
rect 3574 7423 3608 7429
rect 3602 7420 3608 7423
rect 3660 7420 3666 7472
rect 4154 7420 4160 7472
rect 4212 7460 4218 7472
rect 4816 7460 4844 7500
rect 6086 7488 6092 7500
rect 6144 7488 6150 7540
rect 7374 7488 7380 7540
rect 7432 7488 7438 7540
rect 7834 7488 7840 7540
rect 7892 7528 7898 7540
rect 7892 7500 8616 7528
rect 7892 7488 7898 7500
rect 6546 7460 6552 7472
rect 4212 7432 4844 7460
rect 4908 7432 6552 7460
rect 4212 7420 4218 7432
rect 4908 7404 4936 7432
rect 6546 7420 6552 7432
rect 6604 7420 6610 7472
rect 7392 7460 7420 7488
rect 8386 7460 8392 7472
rect 7024 7432 8392 7460
rect 1765 7395 1823 7401
rect 1765 7392 1777 7395
rect 1688 7364 1777 7392
rect 1765 7361 1777 7364
rect 1811 7361 1823 7395
rect 1765 7355 1823 7361
rect 1946 7352 1952 7404
rect 2004 7352 2010 7404
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 4890 7392 4896 7404
rect 2547 7364 4896 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 4982 7352 4988 7404
rect 5040 7352 5046 7404
rect 5902 7352 5908 7404
rect 5960 7401 5966 7404
rect 5960 7355 5972 7401
rect 5960 7352 5966 7355
rect 6270 7352 6276 7404
rect 6328 7352 6334 7404
rect 7024 7401 7052 7432
rect 8386 7420 8392 7432
rect 8444 7420 8450 7472
rect 8588 7460 8616 7500
rect 9858 7488 9864 7540
rect 9916 7488 9922 7540
rect 11330 7528 11336 7540
rect 9968 7500 11336 7528
rect 8726 7463 8784 7469
rect 8726 7460 8738 7463
rect 8588 7432 8738 7460
rect 8726 7429 8738 7432
rect 8772 7429 8784 7463
rect 8726 7423 8784 7429
rect 7009 7395 7067 7401
rect 7009 7361 7021 7395
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 7276 7395 7334 7401
rect 7276 7361 7288 7395
rect 7322 7392 7334 7395
rect 8202 7392 8208 7404
rect 7322 7364 8208 7392
rect 7322 7361 7334 7364
rect 7276 7355 7334 7361
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 9968 7392 9996 7500
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 11440 7500 11744 7528
rect 11440 7460 11468 7500
rect 11348 7432 11468 7460
rect 11348 7401 11376 7432
rect 11514 7420 11520 7472
rect 11572 7420 11578 7472
rect 11716 7460 11744 7500
rect 11790 7488 11796 7540
rect 11848 7528 11854 7540
rect 12069 7531 12127 7537
rect 12069 7528 12081 7531
rect 11848 7500 12081 7528
rect 11848 7488 11854 7500
rect 12069 7497 12081 7500
rect 12115 7497 12127 7531
rect 12069 7491 12127 7497
rect 13538 7488 13544 7540
rect 13596 7488 13602 7540
rect 14274 7488 14280 7540
rect 14332 7528 14338 7540
rect 14737 7531 14795 7537
rect 14737 7528 14749 7531
rect 14332 7500 14749 7528
rect 14332 7488 14338 7500
rect 14737 7497 14749 7500
rect 14783 7497 14795 7531
rect 14737 7491 14795 7497
rect 15562 7488 15568 7540
rect 15620 7528 15626 7540
rect 16301 7531 16359 7537
rect 16301 7528 16313 7531
rect 15620 7500 16313 7528
rect 15620 7488 15626 7500
rect 16301 7497 16313 7500
rect 16347 7497 16359 7531
rect 16301 7491 16359 7497
rect 16758 7488 16764 7540
rect 16816 7528 16822 7540
rect 21082 7528 21088 7540
rect 16816 7500 21088 7528
rect 16816 7488 16822 7500
rect 21082 7488 21088 7500
rect 21140 7488 21146 7540
rect 21266 7488 21272 7540
rect 21324 7488 21330 7540
rect 21450 7488 21456 7540
rect 21508 7488 21514 7540
rect 14461 7463 14519 7469
rect 14461 7460 14473 7463
rect 11716 7432 14473 7460
rect 14461 7429 14473 7432
rect 14507 7429 14519 7463
rect 14461 7423 14519 7429
rect 16132 7432 20668 7460
rect 8352 7364 9996 7392
rect 11077 7395 11135 7401
rect 8352 7352 8358 7364
rect 11077 7361 11089 7395
rect 11123 7392 11135 7395
rect 11333 7395 11391 7401
rect 11123 7364 11284 7392
rect 11123 7361 11135 7364
rect 11077 7355 11135 7361
rect 2685 7327 2743 7333
rect 2685 7293 2697 7327
rect 2731 7324 2743 7327
rect 3050 7324 3056 7336
rect 2731 7296 3056 7324
rect 2731 7293 2743 7296
rect 2685 7287 2743 7293
rect 3050 7284 3056 7296
rect 3108 7284 3114 7336
rect 3142 7284 3148 7336
rect 3200 7324 3206 7336
rect 3329 7327 3387 7333
rect 3329 7324 3341 7327
rect 3200 7296 3341 7324
rect 3200 7284 3206 7296
rect 3329 7293 3341 7296
rect 3375 7293 3387 7327
rect 3329 7287 3387 7293
rect 1673 7259 1731 7265
rect 1673 7225 1685 7259
rect 1719 7256 1731 7259
rect 1719 7228 3372 7256
rect 1719 7225 1731 7228
rect 1673 7219 1731 7225
rect 3344 7188 3372 7228
rect 4430 7216 4436 7268
rect 4488 7216 4494 7268
rect 4801 7259 4859 7265
rect 4801 7225 4813 7259
rect 4847 7256 4859 7259
rect 5000 7256 5028 7352
rect 6181 7327 6239 7333
rect 6181 7293 6193 7327
rect 6227 7324 6239 7327
rect 6288 7324 6316 7352
rect 6227 7296 6316 7324
rect 6227 7293 6239 7296
rect 6181 7287 6239 7293
rect 6822 7284 6828 7336
rect 6880 7324 6886 7336
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 6880 7296 6929 7324
rect 6880 7284 6886 7296
rect 6917 7293 6929 7296
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 8386 7284 8392 7336
rect 8444 7324 8450 7336
rect 8481 7327 8539 7333
rect 8481 7324 8493 7327
rect 8444 7296 8493 7324
rect 8444 7284 8450 7296
rect 8481 7293 8493 7296
rect 8527 7293 8539 7327
rect 11256 7324 11284 7364
rect 11333 7361 11345 7395
rect 11379 7361 11391 7395
rect 11532 7392 11560 7420
rect 11532 7364 11652 7392
rect 11333 7355 11391 7361
rect 11514 7324 11520 7336
rect 11256 7296 11520 7324
rect 8481 7287 8539 7293
rect 11514 7284 11520 7296
rect 11572 7284 11578 7336
rect 11624 7333 11652 7364
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 12417 7395 12475 7401
rect 12417 7392 12429 7395
rect 12124 7364 12429 7392
rect 12124 7352 12130 7364
rect 12417 7361 12429 7364
rect 12463 7361 12475 7395
rect 12417 7355 12475 7361
rect 12710 7352 12716 7404
rect 12768 7392 12774 7404
rect 13633 7395 13691 7401
rect 13633 7392 13645 7395
rect 12768 7364 13645 7392
rect 12768 7352 12774 7364
rect 13633 7361 13645 7364
rect 13679 7361 13691 7395
rect 13633 7355 13691 7361
rect 14366 7352 14372 7404
rect 14424 7352 14430 7404
rect 15838 7352 15844 7404
rect 15896 7401 15902 7404
rect 16132 7401 16160 7432
rect 15896 7355 15908 7401
rect 16117 7395 16175 7401
rect 16117 7361 16129 7395
rect 16163 7361 16175 7395
rect 16117 7355 16175 7361
rect 16209 7395 16267 7401
rect 16209 7361 16221 7395
rect 16255 7392 16267 7395
rect 17793 7395 17851 7401
rect 16255 7364 16344 7392
rect 16255 7361 16267 7364
rect 16209 7355 16267 7361
rect 15896 7352 15902 7355
rect 11609 7327 11667 7333
rect 11609 7293 11621 7327
rect 11655 7324 11667 7327
rect 11790 7324 11796 7336
rect 11655 7296 11796 7324
rect 11655 7293 11667 7296
rect 11609 7287 11667 7293
rect 11790 7284 11796 7296
rect 11848 7284 11854 7336
rect 12161 7327 12219 7333
rect 12161 7293 12173 7327
rect 12207 7293 12219 7327
rect 12161 7287 12219 7293
rect 4847 7228 5028 7256
rect 6641 7259 6699 7265
rect 4847 7225 4859 7228
rect 4801 7219 4859 7225
rect 6641 7225 6653 7259
rect 6687 7225 6699 7259
rect 6641 7219 6699 7225
rect 8220 7228 8524 7256
rect 4448 7188 4476 7216
rect 3344 7160 4476 7188
rect 4614 7148 4620 7200
rect 4672 7188 4678 7200
rect 4709 7191 4767 7197
rect 4709 7188 4721 7191
rect 4672 7160 4721 7188
rect 4672 7148 4678 7160
rect 4709 7157 4721 7160
rect 4755 7157 4767 7191
rect 4709 7151 4767 7157
rect 5534 7148 5540 7200
rect 5592 7188 5598 7200
rect 6457 7191 6515 7197
rect 6457 7188 6469 7191
rect 5592 7160 6469 7188
rect 5592 7148 5598 7160
rect 6457 7157 6469 7160
rect 6503 7157 6515 7191
rect 6656 7188 6684 7219
rect 8220 7200 8248 7228
rect 8110 7188 8116 7200
rect 6656 7160 8116 7188
rect 6457 7151 6515 7157
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 8202 7148 8208 7200
rect 8260 7148 8266 7200
rect 8386 7148 8392 7200
rect 8444 7148 8450 7200
rect 8496 7188 8524 7228
rect 11882 7216 11888 7268
rect 11940 7216 11946 7268
rect 9858 7188 9864 7200
rect 8496 7160 9864 7188
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 9950 7148 9956 7200
rect 10008 7148 10014 7200
rect 12176 7188 12204 7287
rect 13446 7284 13452 7336
rect 13504 7324 13510 7336
rect 14277 7327 14335 7333
rect 14277 7324 14289 7327
rect 13504 7296 14289 7324
rect 13504 7284 13510 7296
rect 14277 7293 14289 7296
rect 14323 7293 14335 7327
rect 14277 7287 14335 7293
rect 13078 7188 13084 7200
rect 12176 7160 13084 7188
rect 13078 7148 13084 7160
rect 13136 7148 13142 7200
rect 13538 7148 13544 7200
rect 13596 7188 13602 7200
rect 16316 7188 16344 7364
rect 17793 7361 17805 7395
rect 17839 7392 17851 7395
rect 17839 7364 18184 7392
rect 17839 7361 17851 7364
rect 17793 7355 17851 7361
rect 18046 7284 18052 7336
rect 18104 7284 18110 7336
rect 18156 7265 18184 7364
rect 18322 7352 18328 7404
rect 18380 7392 18386 7404
rect 19254 7395 19312 7401
rect 19254 7392 19266 7395
rect 18380 7364 19266 7392
rect 18380 7352 18386 7364
rect 19254 7361 19266 7364
rect 19300 7361 19312 7395
rect 19254 7355 19312 7361
rect 19426 7352 19432 7404
rect 19484 7392 19490 7404
rect 19521 7395 19579 7401
rect 19521 7392 19533 7395
rect 19484 7364 19533 7392
rect 19484 7352 19490 7364
rect 19521 7361 19533 7364
rect 19567 7361 19579 7395
rect 19521 7355 19579 7361
rect 19702 7352 19708 7404
rect 19760 7392 19766 7404
rect 19869 7395 19927 7401
rect 19869 7392 19881 7395
rect 19760 7364 19881 7392
rect 19760 7352 19766 7364
rect 19869 7361 19881 7364
rect 19915 7361 19927 7395
rect 19869 7355 19927 7361
rect 19610 7284 19616 7336
rect 19668 7284 19674 7336
rect 20640 7324 20668 7432
rect 21100 7392 21128 7488
rect 21284 7460 21312 7488
rect 21284 7432 21588 7460
rect 21560 7401 21588 7432
rect 23290 7420 23296 7472
rect 23348 7420 23354 7472
rect 21269 7395 21327 7401
rect 21269 7392 21281 7395
rect 21100 7364 21281 7392
rect 21269 7361 21281 7364
rect 21315 7361 21327 7395
rect 21269 7355 21327 7361
rect 21545 7395 21603 7401
rect 21545 7361 21557 7395
rect 21591 7361 21603 7395
rect 21545 7355 21603 7361
rect 21910 7352 21916 7404
rect 21968 7352 21974 7404
rect 22945 7395 23003 7401
rect 22945 7361 22957 7395
rect 22991 7392 23003 7395
rect 23106 7392 23112 7404
rect 22991 7364 23112 7392
rect 22991 7361 23003 7364
rect 22945 7355 23003 7361
rect 23106 7352 23112 7364
rect 23164 7352 23170 7404
rect 23308 7391 23336 7420
rect 23285 7385 23343 7391
rect 21177 7327 21235 7333
rect 21177 7324 21189 7327
rect 20640 7296 21189 7324
rect 21177 7293 21189 7296
rect 21223 7293 21235 7327
rect 21177 7287 21235 7293
rect 18141 7259 18199 7265
rect 18141 7225 18153 7259
rect 18187 7225 18199 7259
rect 18141 7219 18199 7225
rect 20993 7259 21051 7265
rect 20993 7225 21005 7259
rect 21039 7256 21051 7259
rect 21450 7256 21456 7268
rect 21039 7228 21456 7256
rect 21039 7225 21051 7228
rect 20993 7219 21051 7225
rect 21450 7216 21456 7228
rect 21508 7256 21514 7268
rect 21928 7256 21956 7352
rect 23285 7351 23297 7385
rect 23331 7351 23343 7385
rect 23285 7345 23343 7351
rect 23201 7327 23259 7333
rect 23201 7293 23213 7327
rect 23247 7293 23259 7327
rect 23201 7287 23259 7293
rect 21508 7228 21956 7256
rect 23216 7256 23244 7287
rect 23385 7259 23443 7265
rect 23385 7256 23397 7259
rect 23216 7228 23397 7256
rect 21508 7216 21514 7228
rect 23385 7225 23397 7228
rect 23431 7225 23443 7259
rect 23385 7219 23443 7225
rect 13596 7160 16344 7188
rect 16669 7191 16727 7197
rect 13596 7148 13602 7160
rect 16669 7157 16681 7191
rect 16715 7188 16727 7191
rect 16942 7188 16948 7200
rect 16715 7160 16948 7188
rect 16715 7157 16727 7160
rect 16669 7151 16727 7157
rect 16942 7148 16948 7160
rect 17000 7148 17006 7200
rect 21821 7191 21879 7197
rect 21821 7157 21833 7191
rect 21867 7188 21879 7191
rect 23474 7188 23480 7200
rect 21867 7160 23480 7188
rect 21867 7157 21879 7160
rect 21821 7151 21879 7157
rect 23474 7148 23480 7160
rect 23532 7148 23538 7200
rect 1104 7098 23828 7120
rect 1104 7046 1918 7098
rect 1970 7046 1982 7098
rect 2034 7046 2046 7098
rect 2098 7046 2110 7098
rect 2162 7046 2174 7098
rect 2226 7046 2238 7098
rect 2290 7046 7918 7098
rect 7970 7046 7982 7098
rect 8034 7046 8046 7098
rect 8098 7046 8110 7098
rect 8162 7046 8174 7098
rect 8226 7046 8238 7098
rect 8290 7046 13918 7098
rect 13970 7046 13982 7098
rect 14034 7046 14046 7098
rect 14098 7046 14110 7098
rect 14162 7046 14174 7098
rect 14226 7046 14238 7098
rect 14290 7046 19918 7098
rect 19970 7046 19982 7098
rect 20034 7046 20046 7098
rect 20098 7046 20110 7098
rect 20162 7046 20174 7098
rect 20226 7046 20238 7098
rect 20290 7046 23828 7098
rect 1104 7024 23828 7046
rect 1302 6944 1308 6996
rect 1360 6944 1366 6996
rect 1581 6987 1639 6993
rect 1581 6953 1593 6987
rect 1627 6984 1639 6987
rect 1670 6984 1676 6996
rect 1627 6956 1676 6984
rect 1627 6953 1639 6956
rect 1581 6947 1639 6953
rect 1670 6944 1676 6956
rect 1728 6944 1734 6996
rect 1762 6944 1768 6996
rect 1820 6944 1826 6996
rect 2041 6987 2099 6993
rect 2041 6953 2053 6987
rect 2087 6984 2099 6987
rect 2406 6984 2412 6996
rect 2087 6956 2412 6984
rect 2087 6953 2099 6956
rect 2041 6947 2099 6953
rect 2406 6944 2412 6956
rect 2464 6944 2470 6996
rect 3881 6987 3939 6993
rect 3881 6953 3893 6987
rect 3927 6984 3939 6987
rect 4154 6984 4160 6996
rect 3927 6956 4160 6984
rect 3927 6953 3939 6956
rect 3881 6947 3939 6953
rect 4154 6944 4160 6956
rect 4212 6944 4218 6996
rect 4614 6984 4620 6996
rect 4356 6956 4620 6984
rect 1320 6848 1348 6944
rect 1780 6916 1808 6944
rect 1780 6888 1900 6916
rect 1320 6820 1440 6848
rect 1412 6789 1440 6820
rect 1486 6808 1492 6860
rect 1544 6848 1550 6860
rect 1765 6851 1823 6857
rect 1765 6848 1777 6851
rect 1544 6820 1777 6848
rect 1544 6808 1550 6820
rect 1765 6817 1777 6820
rect 1811 6817 1823 6851
rect 1765 6811 1823 6817
rect 1872 6789 1900 6888
rect 3050 6876 3056 6928
rect 3108 6876 3114 6928
rect 4356 6916 4384 6956
rect 4614 6944 4620 6956
rect 4672 6944 4678 6996
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 10502 6984 10508 6996
rect 8444 6956 10508 6984
rect 8444 6944 8450 6956
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 15473 6987 15531 6993
rect 15473 6953 15485 6987
rect 15519 6984 15531 6987
rect 16298 6984 16304 6996
rect 15519 6956 16304 6984
rect 15519 6953 15531 6956
rect 15473 6947 15531 6953
rect 16298 6944 16304 6956
rect 16356 6944 16362 6996
rect 18785 6987 18843 6993
rect 18785 6953 18797 6987
rect 18831 6984 18843 6987
rect 18874 6984 18880 6996
rect 18831 6956 18880 6984
rect 18831 6953 18843 6956
rect 18785 6947 18843 6953
rect 18874 6944 18880 6956
rect 18932 6944 18938 6996
rect 19426 6984 19432 6996
rect 19260 6956 19432 6984
rect 4080 6888 4384 6916
rect 2774 6808 2780 6860
rect 2832 6808 2838 6860
rect 2961 6851 3019 6857
rect 2961 6817 2973 6851
rect 3007 6848 3019 6851
rect 3068 6848 3096 6876
rect 3007 6820 3096 6848
rect 3007 6817 3019 6820
rect 2961 6811 3019 6817
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6749 1915 6783
rect 1857 6743 1915 6749
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6780 2007 6783
rect 2498 6780 2504 6792
rect 1995 6752 2504 6780
rect 1995 6749 2007 6752
rect 1949 6743 2007 6749
rect 2498 6740 2504 6752
rect 2556 6740 2562 6792
rect 2593 6783 2651 6789
rect 2593 6749 2605 6783
rect 2639 6749 2651 6783
rect 2593 6743 2651 6749
rect 2608 6712 2636 6743
rect 2866 6740 2872 6792
rect 2924 6740 2930 6792
rect 3786 6780 3792 6792
rect 2976 6752 3792 6780
rect 2976 6712 3004 6752
rect 3786 6740 3792 6752
rect 3844 6740 3850 6792
rect 4080 6789 4108 6888
rect 8294 6876 8300 6928
rect 8352 6916 8358 6928
rect 9033 6919 9091 6925
rect 9033 6916 9045 6919
rect 8352 6888 9045 6916
rect 8352 6876 8358 6888
rect 9033 6885 9045 6888
rect 9079 6885 9091 6919
rect 9033 6879 9091 6885
rect 9217 6919 9275 6925
rect 9217 6885 9229 6919
rect 9263 6916 9275 6919
rect 9398 6916 9404 6928
rect 9263 6888 9404 6916
rect 9263 6885 9275 6888
rect 9217 6879 9275 6885
rect 9398 6876 9404 6888
rect 9456 6876 9462 6928
rect 4157 6851 4215 6857
rect 4157 6817 4169 6851
rect 4203 6848 4215 6851
rect 4246 6848 4252 6860
rect 4203 6820 4252 6848
rect 4203 6817 4215 6820
rect 4157 6811 4215 6817
rect 4246 6808 4252 6820
rect 4304 6808 4310 6860
rect 8478 6808 8484 6860
rect 8536 6848 8542 6860
rect 9490 6848 9496 6860
rect 8536 6820 9496 6848
rect 8536 6808 8542 6820
rect 9490 6808 9496 6820
rect 9548 6848 9554 6860
rect 9585 6851 9643 6857
rect 9585 6848 9597 6851
rect 9548 6820 9597 6848
rect 9548 6808 9554 6820
rect 9585 6817 9597 6820
rect 9631 6817 9643 6851
rect 19260 6848 19288 6956
rect 19426 6944 19432 6956
rect 19484 6944 19490 6996
rect 22002 6944 22008 6996
rect 22060 6984 22066 6996
rect 22278 6984 22284 6996
rect 22060 6956 22284 6984
rect 22060 6944 22066 6956
rect 22278 6944 22284 6956
rect 22336 6944 22342 6996
rect 22186 6848 22192 6860
rect 9585 6811 9643 6817
rect 18800 6820 19288 6848
rect 21928 6820 22192 6848
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6780 4399 6783
rect 5810 6780 5816 6792
rect 4387 6752 5816 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 7282 6740 7288 6792
rect 7340 6740 7346 6792
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6780 11115 6783
rect 12434 6780 12440 6792
rect 11103 6752 12440 6780
rect 11103 6749 11115 6752
rect 11057 6743 11115 6749
rect 12434 6740 12440 6752
rect 12492 6740 12498 6792
rect 13814 6740 13820 6792
rect 13872 6780 13878 6792
rect 14090 6780 14096 6792
rect 13872 6752 14096 6780
rect 13872 6740 13878 6752
rect 14090 6740 14096 6752
rect 14148 6740 14154 6792
rect 14366 6789 14372 6792
rect 14360 6780 14372 6789
rect 14327 6752 14372 6780
rect 14360 6743 14372 6752
rect 14366 6740 14372 6743
rect 14424 6740 14430 6792
rect 16945 6783 17003 6789
rect 16945 6749 16957 6783
rect 16991 6780 17003 6783
rect 17221 6783 17279 6789
rect 17221 6780 17233 6783
rect 16991 6752 17233 6780
rect 16991 6749 17003 6752
rect 16945 6743 17003 6749
rect 17221 6749 17233 6752
rect 17267 6780 17279 6783
rect 18800 6780 18828 6820
rect 17267 6752 18828 6780
rect 18877 6783 18935 6789
rect 17267 6749 17279 6752
rect 17221 6743 17279 6749
rect 18877 6749 18889 6783
rect 18923 6780 18935 6783
rect 18966 6780 18972 6792
rect 18923 6752 18972 6780
rect 18923 6749 18935 6752
rect 18877 6743 18935 6749
rect 18966 6740 18972 6752
rect 19024 6740 19030 6792
rect 19242 6740 19248 6792
rect 19300 6740 19306 6792
rect 20717 6783 20775 6789
rect 20717 6749 20729 6783
rect 20763 6780 20775 6783
rect 21358 6780 21364 6792
rect 20763 6752 21364 6780
rect 20763 6749 20775 6752
rect 20717 6743 20775 6749
rect 21358 6740 21364 6752
rect 21416 6740 21422 6792
rect 4586 6715 4644 6721
rect 4586 6712 4598 6715
rect 2608 6684 3004 6712
rect 3804 6684 4598 6712
rect 2501 6647 2559 6653
rect 2501 6613 2513 6647
rect 2547 6644 2559 6647
rect 2682 6644 2688 6656
rect 2547 6616 2688 6644
rect 2547 6613 2559 6616
rect 2501 6607 2559 6613
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 3605 6647 3663 6653
rect 3605 6613 3617 6647
rect 3651 6644 3663 6647
rect 3804 6644 3832 6684
rect 4586 6681 4598 6684
rect 4632 6681 4644 6715
rect 4586 6675 4644 6681
rect 7552 6715 7610 6721
rect 7552 6681 7564 6715
rect 7598 6712 7610 6715
rect 7650 6712 7656 6724
rect 7598 6684 7656 6712
rect 7598 6681 7610 6684
rect 7552 6675 7610 6681
rect 7650 6672 7656 6684
rect 7708 6672 7714 6724
rect 9493 6715 9551 6721
rect 9493 6712 9505 6715
rect 8404 6684 9505 6712
rect 3651 6616 3832 6644
rect 5721 6647 5779 6653
rect 3651 6613 3663 6616
rect 3605 6607 3663 6613
rect 5721 6613 5733 6647
rect 5767 6644 5779 6647
rect 6270 6644 6276 6656
rect 5767 6616 6276 6644
rect 5767 6613 5779 6616
rect 5721 6607 5779 6613
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 6822 6604 6828 6656
rect 6880 6644 6886 6656
rect 8404 6644 8432 6684
rect 9493 6681 9505 6684
rect 9539 6712 9551 6715
rect 9674 6712 9680 6724
rect 9539 6684 9680 6712
rect 9539 6681 9551 6684
rect 9493 6675 9551 6681
rect 9674 6672 9680 6684
rect 9732 6672 9738 6724
rect 9852 6715 9910 6721
rect 9852 6681 9864 6715
rect 9898 6712 9910 6715
rect 9950 6712 9956 6724
rect 9898 6684 9956 6712
rect 9898 6681 9910 6684
rect 9852 6675 9910 6681
rect 9950 6672 9956 6684
rect 10008 6672 10014 6724
rect 11324 6715 11382 6721
rect 11324 6681 11336 6715
rect 11370 6681 11382 6715
rect 11324 6675 11382 6681
rect 16700 6715 16758 6721
rect 16700 6681 16712 6715
rect 16746 6712 16758 6715
rect 17488 6715 17546 6721
rect 16746 6684 17448 6712
rect 16746 6681 16758 6684
rect 16700 6675 16758 6681
rect 6880 6616 8432 6644
rect 6880 6604 6886 6616
rect 8478 6604 8484 6656
rect 8536 6644 8542 6656
rect 8665 6647 8723 6653
rect 8665 6644 8677 6647
rect 8536 6616 8677 6644
rect 8536 6604 8542 6616
rect 8665 6613 8677 6616
rect 8711 6613 8723 6647
rect 8665 6607 8723 6613
rect 10965 6647 11023 6653
rect 10965 6613 10977 6647
rect 11011 6644 11023 6647
rect 11054 6644 11060 6656
rect 11011 6616 11060 6644
rect 11011 6613 11023 6616
rect 10965 6607 11023 6613
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 11348 6644 11376 6675
rect 11296 6616 11376 6644
rect 12437 6647 12495 6653
rect 11296 6604 11302 6616
rect 12437 6613 12449 6647
rect 12483 6644 12495 6647
rect 13354 6644 13360 6656
rect 12483 6616 13360 6644
rect 12483 6613 12495 6616
rect 12437 6607 12495 6613
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 15565 6647 15623 6653
rect 15565 6613 15577 6647
rect 15611 6644 15623 6647
rect 15746 6644 15752 6656
rect 15611 6616 15752 6644
rect 15611 6613 15623 6616
rect 15565 6607 15623 6613
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 17420 6644 17448 6684
rect 17488 6681 17500 6715
rect 17534 6712 17546 6715
rect 17862 6712 17868 6724
rect 17534 6684 17868 6712
rect 17534 6681 17546 6684
rect 17488 6675 17546 6681
rect 17862 6672 17868 6684
rect 17920 6672 17926 6724
rect 19518 6721 19524 6724
rect 19512 6675 19524 6721
rect 19518 6672 19524 6675
rect 19576 6672 19582 6724
rect 19702 6672 19708 6724
rect 19760 6672 19766 6724
rect 20984 6715 21042 6721
rect 20984 6681 20996 6715
rect 21030 6712 21042 6715
rect 21928 6712 21956 6820
rect 22186 6808 22192 6820
rect 22244 6808 22250 6860
rect 22922 6808 22928 6860
rect 22980 6848 22986 6860
rect 23109 6851 23167 6857
rect 23109 6848 23121 6851
rect 22980 6820 23121 6848
rect 22980 6808 22986 6820
rect 23109 6817 23121 6820
rect 23155 6817 23167 6851
rect 23109 6811 23167 6817
rect 22833 6783 22891 6789
rect 22833 6780 22845 6783
rect 21030 6684 21956 6712
rect 22020 6752 22845 6780
rect 21030 6681 21042 6684
rect 20984 6675 21042 6681
rect 17678 6644 17684 6656
rect 17420 6616 17684 6644
rect 17678 6604 17684 6616
rect 17736 6604 17742 6656
rect 18601 6647 18659 6653
rect 18601 6613 18613 6647
rect 18647 6644 18659 6647
rect 19720 6644 19748 6672
rect 18647 6616 19748 6644
rect 20625 6647 20683 6653
rect 18647 6613 18659 6616
rect 18601 6607 18659 6613
rect 20625 6613 20637 6647
rect 20671 6644 20683 6647
rect 22020 6644 22048 6752
rect 22833 6749 22845 6752
rect 22879 6749 22891 6783
rect 22833 6743 22891 6749
rect 20671 6616 22048 6644
rect 22097 6647 22155 6653
rect 20671 6613 20683 6616
rect 20625 6607 20683 6613
rect 22097 6613 22109 6647
rect 22143 6644 22155 6647
rect 22554 6644 22560 6656
rect 22143 6616 22560 6644
rect 22143 6613 22155 6616
rect 22097 6607 22155 6613
rect 22554 6604 22560 6616
rect 22612 6604 22618 6656
rect 1104 6554 23828 6576
rect 1104 6502 2658 6554
rect 2710 6502 2722 6554
rect 2774 6502 2786 6554
rect 2838 6502 2850 6554
rect 2902 6502 2914 6554
rect 2966 6502 2978 6554
rect 3030 6502 8658 6554
rect 8710 6502 8722 6554
rect 8774 6502 8786 6554
rect 8838 6502 8850 6554
rect 8902 6502 8914 6554
rect 8966 6502 8978 6554
rect 9030 6502 14658 6554
rect 14710 6502 14722 6554
rect 14774 6502 14786 6554
rect 14838 6502 14850 6554
rect 14902 6502 14914 6554
rect 14966 6502 14978 6554
rect 15030 6502 20658 6554
rect 20710 6502 20722 6554
rect 20774 6502 20786 6554
rect 20838 6502 20850 6554
rect 20902 6502 20914 6554
rect 20966 6502 20978 6554
rect 21030 6502 23828 6554
rect 1104 6480 23828 6502
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 1673 6443 1731 6449
rect 1673 6440 1685 6443
rect 1452 6412 1685 6440
rect 1452 6400 1458 6412
rect 1673 6409 1685 6412
rect 1719 6409 1731 6443
rect 4709 6443 4767 6449
rect 1673 6403 1731 6409
rect 3600 6412 4660 6440
rect 1578 6332 1584 6384
rect 1636 6332 1642 6384
rect 3600 6372 3628 6412
rect 4522 6372 4528 6384
rect 3344 6344 3628 6372
rect 3804 6344 4528 6372
rect 1596 6304 1624 6332
rect 3344 6313 3372 6344
rect 1765 6307 1823 6313
rect 1765 6304 1777 6307
rect 1596 6276 1777 6304
rect 1765 6273 1777 6276
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 2124 6307 2182 6313
rect 2124 6273 2136 6307
rect 2170 6304 2182 6307
rect 3329 6307 3387 6313
rect 2170 6276 3096 6304
rect 2170 6273 2182 6276
rect 2124 6267 2182 6273
rect 3068 6248 3096 6276
rect 3329 6273 3341 6307
rect 3375 6273 3387 6307
rect 3329 6267 3387 6273
rect 3596 6307 3654 6313
rect 3596 6273 3608 6307
rect 3642 6304 3654 6307
rect 3804 6304 3832 6344
rect 4522 6332 4528 6344
rect 4580 6332 4586 6384
rect 4632 6372 4660 6412
rect 4709 6409 4721 6443
rect 4755 6440 4767 6443
rect 4755 6412 4844 6440
rect 4755 6409 4767 6412
rect 4709 6403 4767 6409
rect 4632 6344 4752 6372
rect 4724 6316 4752 6344
rect 3642 6276 3832 6304
rect 3642 6273 3654 6276
rect 3596 6267 3654 6273
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6205 1915 6239
rect 1857 6199 1915 6205
rect 1872 6100 1900 6199
rect 3050 6196 3056 6248
rect 3108 6196 3114 6248
rect 3344 6168 3372 6267
rect 4338 6264 4344 6316
rect 4396 6304 4402 6316
rect 4614 6304 4620 6316
rect 4396 6276 4620 6304
rect 4396 6264 4402 6276
rect 4614 6264 4620 6276
rect 4672 6264 4678 6316
rect 4706 6264 4712 6316
rect 4764 6264 4770 6316
rect 4816 6304 4844 6412
rect 6178 6400 6184 6452
rect 6236 6440 6242 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 6236 6412 6561 6440
rect 6236 6400 6242 6412
rect 6549 6409 6561 6412
rect 6595 6409 6607 6443
rect 6549 6403 6607 6409
rect 6638 6400 6644 6452
rect 6696 6440 6702 6452
rect 6825 6443 6883 6449
rect 6825 6440 6837 6443
rect 6696 6412 6837 6440
rect 6696 6400 6702 6412
rect 6825 6409 6837 6412
rect 6871 6409 6883 6443
rect 6825 6403 6883 6409
rect 6914 6400 6920 6452
rect 6972 6400 6978 6452
rect 7006 6400 7012 6452
rect 7064 6400 7070 6452
rect 9858 6400 9864 6452
rect 9916 6400 9922 6452
rect 10318 6400 10324 6452
rect 10376 6400 10382 6452
rect 11330 6400 11336 6452
rect 11388 6440 11394 6452
rect 11517 6443 11575 6449
rect 11517 6440 11529 6443
rect 11388 6412 11529 6440
rect 11388 6400 11394 6412
rect 11517 6409 11529 6412
rect 11563 6409 11575 6443
rect 11517 6403 11575 6409
rect 12529 6443 12587 6449
rect 12529 6409 12541 6443
rect 12575 6409 12587 6443
rect 12529 6403 12587 6409
rect 6932 6372 6960 6400
rect 6656 6344 6960 6372
rect 6656 6313 6684 6344
rect 5057 6307 5115 6313
rect 5057 6304 5069 6307
rect 4816 6276 5069 6304
rect 5057 6273 5069 6276
rect 5103 6273 5115 6307
rect 5057 6267 5115 6273
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6304 6975 6307
rect 7024 6304 7052 6400
rect 6963 6276 7052 6304
rect 6963 6273 6975 6276
rect 6917 6267 6975 6273
rect 7098 6264 7104 6316
rect 7156 6304 7162 6316
rect 7265 6307 7323 6313
rect 7265 6304 7277 6307
rect 7156 6276 7277 6304
rect 7156 6264 7162 6276
rect 7265 6273 7277 6276
rect 7311 6273 7323 6307
rect 7265 6267 7323 6273
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 7616 6276 8493 6304
rect 7616 6264 7622 6276
rect 8481 6273 8493 6276
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 8748 6307 8806 6313
rect 8748 6273 8760 6307
rect 8794 6304 8806 6307
rect 9030 6304 9036 6316
rect 8794 6276 9036 6304
rect 8794 6273 8806 6276
rect 8748 6267 8806 6273
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 9490 6264 9496 6316
rect 9548 6304 9554 6316
rect 9950 6304 9956 6316
rect 9548 6276 9956 6304
rect 9548 6264 9554 6276
rect 9950 6264 9956 6276
rect 10008 6264 10014 6316
rect 10226 6313 10232 6316
rect 10220 6304 10232 6313
rect 10187 6276 10232 6304
rect 10220 6267 10232 6276
rect 10226 6264 10232 6267
rect 10284 6264 10290 6316
rect 10336 6304 10364 6400
rect 12544 6372 12572 6403
rect 13630 6400 13636 6452
rect 13688 6440 13694 6452
rect 15286 6440 15292 6452
rect 13688 6412 15292 6440
rect 13688 6400 13694 6412
rect 15286 6400 15292 6412
rect 15344 6400 15350 6452
rect 15930 6400 15936 6452
rect 15988 6440 15994 6452
rect 16393 6443 16451 6449
rect 16393 6440 16405 6443
rect 15988 6412 16405 6440
rect 15988 6400 15994 6412
rect 16393 6409 16405 6412
rect 16439 6409 16451 6443
rect 16393 6403 16451 6409
rect 16574 6400 16580 6452
rect 16632 6440 16638 6452
rect 16761 6443 16819 6449
rect 16761 6440 16773 6443
rect 16632 6412 16773 6440
rect 16632 6400 16638 6412
rect 16761 6409 16773 6412
rect 16807 6409 16819 6443
rect 16761 6403 16819 6409
rect 18506 6400 18512 6452
rect 18564 6400 18570 6452
rect 18782 6400 18788 6452
rect 18840 6400 18846 6452
rect 19242 6400 19248 6452
rect 19300 6440 19306 6452
rect 21269 6443 21327 6449
rect 21269 6440 21281 6443
rect 19300 6412 21281 6440
rect 19300 6400 19306 6412
rect 21269 6409 21281 6412
rect 21315 6409 21327 6443
rect 21269 6403 21327 6409
rect 23014 6400 23020 6452
rect 23072 6440 23078 6452
rect 23385 6443 23443 6449
rect 23385 6440 23397 6443
rect 23072 6412 23397 6440
rect 23072 6400 23078 6412
rect 23385 6409 23397 6412
rect 23431 6409 23443 6443
rect 23385 6403 23443 6409
rect 14338 6375 14396 6381
rect 14338 6372 14350 6375
rect 12544 6344 14350 6372
rect 14338 6341 14350 6344
rect 14384 6341 14396 6375
rect 14338 6335 14396 6341
rect 16666 6332 16672 6384
rect 16724 6372 16730 6384
rect 16724 6344 16896 6372
rect 16724 6332 16730 6344
rect 12069 6307 12127 6313
rect 12069 6304 12081 6307
rect 10336 6276 12081 6304
rect 12069 6273 12081 6276
rect 12115 6273 12127 6307
rect 12069 6267 12127 6273
rect 13630 6264 13636 6316
rect 13688 6313 13694 6316
rect 13688 6267 13700 6313
rect 13688 6264 13694 6267
rect 13814 6264 13820 6316
rect 13872 6304 13878 6316
rect 13909 6307 13967 6313
rect 13909 6304 13921 6307
rect 13872 6276 13921 6304
rect 13872 6264 13878 6276
rect 13909 6273 13921 6276
rect 13955 6273 13967 6307
rect 13909 6267 13967 6273
rect 16114 6264 16120 6316
rect 16172 6264 16178 6316
rect 16485 6307 16543 6313
rect 16485 6273 16497 6307
rect 16531 6304 16543 6307
rect 16758 6304 16764 6316
rect 16531 6276 16764 6304
rect 16531 6273 16543 6276
rect 16485 6267 16543 6273
rect 16758 6264 16764 6276
rect 16816 6264 16822 6316
rect 16868 6313 16896 6344
rect 16853 6307 16911 6313
rect 16853 6273 16865 6307
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 18138 6264 18144 6316
rect 18196 6313 18202 6316
rect 18196 6267 18208 6313
rect 18693 6307 18751 6313
rect 18693 6273 18705 6307
rect 18739 6304 18751 6307
rect 18800 6304 18828 6400
rect 20104 6375 20162 6381
rect 20104 6341 20116 6375
rect 20150 6372 20162 6375
rect 20990 6372 20996 6384
rect 20150 6344 20996 6372
rect 20150 6341 20162 6344
rect 20104 6335 20162 6341
rect 20990 6332 20996 6344
rect 21048 6332 21054 6384
rect 18739 6276 18828 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 18196 6264 18202 6267
rect 19794 6264 19800 6316
rect 19852 6304 19858 6316
rect 20441 6307 20499 6313
rect 20441 6304 20453 6307
rect 19852 6276 20453 6304
rect 19852 6264 19858 6276
rect 20441 6273 20453 6276
rect 20487 6273 20499 6307
rect 20441 6267 20499 6273
rect 21085 6307 21143 6313
rect 21085 6273 21097 6307
rect 21131 6304 21143 6307
rect 21174 6304 21180 6316
rect 21131 6276 21180 6304
rect 21131 6273 21143 6276
rect 21085 6267 21143 6273
rect 21174 6264 21180 6276
rect 21232 6264 21238 6316
rect 21266 6264 21272 6316
rect 21324 6304 21330 6316
rect 21361 6307 21419 6313
rect 21361 6304 21373 6307
rect 21324 6276 21373 6304
rect 21324 6264 21330 6276
rect 21361 6273 21373 6276
rect 21407 6304 21419 6307
rect 21637 6307 21695 6313
rect 21637 6304 21649 6307
rect 21407 6276 21649 6304
rect 21407 6273 21419 6276
rect 21361 6267 21419 6273
rect 21637 6273 21649 6276
rect 21683 6273 21695 6307
rect 21637 6267 21695 6273
rect 22945 6307 23003 6313
rect 22945 6273 22957 6307
rect 22991 6304 23003 6307
rect 23106 6304 23112 6316
rect 22991 6276 23112 6304
rect 22991 6273 23003 6276
rect 22945 6267 23003 6273
rect 23106 6264 23112 6276
rect 23164 6264 23170 6316
rect 23293 6307 23351 6313
rect 23293 6273 23305 6307
rect 23339 6304 23351 6307
rect 23382 6304 23388 6316
rect 23339 6276 23388 6304
rect 23339 6273 23351 6276
rect 23293 6267 23351 6273
rect 23382 6264 23388 6276
rect 23440 6264 23446 6316
rect 4801 6239 4859 6245
rect 4801 6205 4813 6239
rect 4847 6205 4859 6239
rect 4801 6199 4859 6205
rect 3160 6140 3372 6168
rect 3160 6100 3188 6140
rect 4338 6128 4344 6180
rect 4396 6168 4402 6180
rect 4816 6168 4844 6199
rect 6546 6196 6552 6248
rect 6604 6236 6610 6248
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 6604 6208 7021 6236
rect 6604 6196 6610 6208
rect 7009 6205 7021 6208
rect 7055 6205 7067 6239
rect 7009 6199 7067 6205
rect 11698 6196 11704 6248
rect 11756 6196 11762 6248
rect 14090 6196 14096 6248
rect 14148 6196 14154 6248
rect 18414 6196 18420 6248
rect 18472 6196 18478 6248
rect 20349 6239 20407 6245
rect 20349 6205 20361 6239
rect 20395 6205 20407 6239
rect 20349 6199 20407 6205
rect 11716 6168 11744 6196
rect 4396 6140 4844 6168
rect 10888 6140 11744 6168
rect 4396 6128 4402 6140
rect 1872 6072 3188 6100
rect 3237 6103 3295 6109
rect 3237 6069 3249 6103
rect 3283 6100 3295 6103
rect 4430 6100 4436 6112
rect 3283 6072 4436 6100
rect 3283 6069 3295 6072
rect 3237 6063 3295 6069
rect 4430 6060 4436 6072
rect 4488 6060 4494 6112
rect 6181 6103 6239 6109
rect 6181 6069 6193 6103
rect 6227 6100 6239 6103
rect 6638 6100 6644 6112
rect 6227 6072 6644 6100
rect 6227 6069 6239 6072
rect 6181 6063 6239 6069
rect 6638 6060 6644 6072
rect 6696 6060 6702 6112
rect 8389 6103 8447 6109
rect 8389 6069 8401 6103
rect 8435 6100 8447 6103
rect 10888 6100 10916 6140
rect 8435 6072 10916 6100
rect 8435 6069 8447 6072
rect 8389 6063 8447 6069
rect 11330 6060 11336 6112
rect 11388 6060 11394 6112
rect 14108 6100 14136 6196
rect 20364 6168 20392 6199
rect 23198 6196 23204 6248
rect 23256 6196 23262 6248
rect 21545 6171 21603 6177
rect 21545 6168 21557 6171
rect 20364 6140 21557 6168
rect 21545 6137 21557 6140
rect 21591 6137 21603 6171
rect 21545 6131 21603 6137
rect 14366 6100 14372 6112
rect 14108 6072 14372 6100
rect 14366 6060 14372 6072
rect 14424 6060 14430 6112
rect 15470 6060 15476 6112
rect 15528 6060 15534 6112
rect 15565 6103 15623 6109
rect 15565 6069 15577 6103
rect 15611 6100 15623 6103
rect 15654 6100 15660 6112
rect 15611 6072 15660 6100
rect 15611 6069 15623 6072
rect 15565 6063 15623 6069
rect 15654 6060 15660 6072
rect 15712 6060 15718 6112
rect 17034 6060 17040 6112
rect 17092 6060 17098 6112
rect 18969 6103 19027 6109
rect 18969 6069 18981 6103
rect 19015 6100 19027 6103
rect 20346 6100 20352 6112
rect 19015 6072 20352 6100
rect 19015 6069 19027 6072
rect 18969 6063 19027 6069
rect 20346 6060 20352 6072
rect 20404 6060 20410 6112
rect 20898 6060 20904 6112
rect 20956 6100 20962 6112
rect 21821 6103 21879 6109
rect 21821 6100 21833 6103
rect 20956 6072 21833 6100
rect 20956 6060 20962 6072
rect 21821 6069 21833 6072
rect 21867 6069 21879 6103
rect 21821 6063 21879 6069
rect 1104 6010 23828 6032
rect 1104 5958 1918 6010
rect 1970 5958 1982 6010
rect 2034 5958 2046 6010
rect 2098 5958 2110 6010
rect 2162 5958 2174 6010
rect 2226 5958 2238 6010
rect 2290 5958 7918 6010
rect 7970 5958 7982 6010
rect 8034 5958 8046 6010
rect 8098 5958 8110 6010
rect 8162 5958 8174 6010
rect 8226 5958 8238 6010
rect 8290 5958 13918 6010
rect 13970 5958 13982 6010
rect 14034 5958 14046 6010
rect 14098 5958 14110 6010
rect 14162 5958 14174 6010
rect 14226 5958 14238 6010
rect 14290 5958 19918 6010
rect 19970 5958 19982 6010
rect 20034 5958 20046 6010
rect 20098 5958 20110 6010
rect 20162 5958 20174 6010
rect 20226 5958 20238 6010
rect 20290 5958 23828 6010
rect 1104 5936 23828 5958
rect 1578 5856 1584 5908
rect 1636 5856 1642 5908
rect 2317 5899 2375 5905
rect 2317 5865 2329 5899
rect 2363 5896 2375 5899
rect 2774 5896 2780 5908
rect 2363 5868 2780 5896
rect 2363 5865 2375 5868
rect 2317 5859 2375 5865
rect 2774 5856 2780 5868
rect 2832 5856 2838 5908
rect 2869 5899 2927 5905
rect 2869 5865 2881 5899
rect 2915 5896 2927 5899
rect 3326 5896 3332 5908
rect 2915 5868 3332 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 3326 5856 3332 5868
rect 3384 5856 3390 5908
rect 3881 5899 3939 5905
rect 3881 5865 3893 5899
rect 3927 5896 3939 5899
rect 4062 5896 4068 5908
rect 3927 5868 4068 5896
rect 3927 5865 3939 5868
rect 3881 5859 3939 5865
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 4157 5899 4215 5905
rect 4157 5865 4169 5899
rect 4203 5896 4215 5899
rect 4246 5896 4252 5908
rect 4203 5868 4252 5896
rect 4203 5865 4215 5868
rect 4157 5859 4215 5865
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 9033 5899 9091 5905
rect 7392 5868 8708 5896
rect 1596 5760 1624 5856
rect 2498 5788 2504 5840
rect 2556 5788 2562 5840
rect 2593 5831 2651 5837
rect 2593 5797 2605 5831
rect 2639 5828 2651 5831
rect 3234 5828 3240 5840
rect 2639 5800 3240 5828
rect 2639 5797 2651 5800
rect 2593 5791 2651 5797
rect 3234 5788 3240 5800
rect 3292 5788 3298 5840
rect 3786 5788 3792 5840
rect 3844 5828 3850 5840
rect 3844 5800 4200 5828
rect 3844 5788 3850 5800
rect 1946 5760 1952 5772
rect 1596 5732 1952 5760
rect 1210 5652 1216 5704
rect 1268 5652 1274 5704
rect 1872 5701 1900 5732
rect 1946 5720 1952 5732
rect 2004 5760 2010 5772
rect 2516 5760 2544 5788
rect 4172 5760 4200 5800
rect 7392 5760 7420 5868
rect 2004 5732 2268 5760
rect 2516 5732 3464 5760
rect 4172 5732 4292 5760
rect 2004 5720 2010 5732
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 1228 5556 1256 5652
rect 1596 5624 1624 5655
rect 2130 5652 2136 5704
rect 2188 5652 2194 5704
rect 2240 5692 2268 5732
rect 2792 5701 2820 5732
rect 2501 5695 2559 5701
rect 2501 5692 2513 5695
rect 2240 5664 2513 5692
rect 2501 5661 2513 5664
rect 2547 5661 2559 5695
rect 2501 5655 2559 5661
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 3050 5652 3056 5704
rect 3108 5692 3114 5704
rect 3436 5701 3464 5732
rect 3237 5695 3295 5701
rect 3237 5692 3249 5695
rect 3108 5664 3249 5692
rect 3108 5652 3114 5664
rect 3237 5661 3249 5664
rect 3283 5661 3295 5695
rect 3237 5655 3295 5661
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5661 3479 5695
rect 3421 5655 3479 5661
rect 3970 5652 3976 5704
rect 4028 5652 4034 5704
rect 4089 5697 4147 5703
rect 4089 5663 4101 5697
rect 4135 5694 4147 5697
rect 4264 5694 4292 5732
rect 7116 5732 7420 5760
rect 8680 5760 8708 5868
rect 9033 5865 9045 5899
rect 9079 5896 9091 5899
rect 9122 5896 9128 5908
rect 9079 5868 9128 5896
rect 9079 5865 9091 5868
rect 9033 5859 9091 5865
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 10318 5896 10324 5908
rect 9324 5868 10324 5896
rect 8757 5831 8815 5837
rect 8757 5797 8769 5831
rect 8803 5828 8815 5831
rect 9324 5828 9352 5868
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 10704 5868 12434 5896
rect 10704 5837 10732 5868
rect 8803 5800 9352 5828
rect 10689 5831 10747 5837
rect 8803 5797 8815 5800
rect 8757 5791 8815 5797
rect 10689 5797 10701 5831
rect 10735 5797 10747 5831
rect 10689 5791 10747 5797
rect 12161 5831 12219 5837
rect 12161 5797 12173 5831
rect 12207 5797 12219 5831
rect 12406 5828 12434 5868
rect 12710 5856 12716 5908
rect 12768 5856 12774 5908
rect 12986 5856 12992 5908
rect 13044 5896 13050 5908
rect 14645 5899 14703 5905
rect 14645 5896 14657 5899
rect 13044 5868 14657 5896
rect 13044 5856 13050 5868
rect 14645 5865 14657 5868
rect 14691 5865 14703 5899
rect 15654 5896 15660 5908
rect 14645 5859 14703 5865
rect 14844 5868 15660 5896
rect 12618 5828 12624 5840
rect 12406 5800 12624 5828
rect 12161 5791 12219 5797
rect 12176 5760 12204 5791
rect 12618 5788 12624 5800
rect 12676 5788 12682 5840
rect 12728 5760 12756 5856
rect 13722 5788 13728 5840
rect 13780 5828 13786 5840
rect 14093 5831 14151 5837
rect 14093 5828 14105 5831
rect 13780 5800 14105 5828
rect 13780 5788 13786 5800
rect 14093 5797 14105 5800
rect 14139 5797 14151 5831
rect 14093 5791 14151 5797
rect 14277 5831 14335 5837
rect 14277 5797 14289 5831
rect 14323 5828 14335 5831
rect 14844 5828 14872 5868
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 18046 5856 18052 5908
rect 18104 5896 18110 5908
rect 18969 5899 19027 5905
rect 18969 5896 18981 5899
rect 18104 5868 18981 5896
rect 18104 5856 18110 5868
rect 18969 5865 18981 5868
rect 19015 5865 19027 5899
rect 18969 5859 19027 5865
rect 19337 5899 19395 5905
rect 19337 5865 19349 5899
rect 19383 5896 19395 5899
rect 19610 5896 19616 5908
rect 19383 5868 19616 5896
rect 19383 5865 19395 5868
rect 19337 5859 19395 5865
rect 19610 5856 19616 5868
rect 19668 5856 19674 5908
rect 20346 5856 20352 5908
rect 20404 5856 20410 5908
rect 20898 5856 20904 5908
rect 20956 5856 20962 5908
rect 20990 5856 20996 5908
rect 21048 5856 21054 5908
rect 21542 5856 21548 5908
rect 21600 5896 21606 5908
rect 21821 5899 21879 5905
rect 21821 5896 21833 5899
rect 21600 5868 21833 5896
rect 21600 5856 21606 5868
rect 21821 5865 21833 5868
rect 21867 5865 21879 5899
rect 21821 5859 21879 5865
rect 22002 5856 22008 5908
rect 22060 5856 22066 5908
rect 14323 5800 14872 5828
rect 14323 5797 14335 5800
rect 14277 5791 14335 5797
rect 18138 5788 18144 5840
rect 18196 5788 18202 5840
rect 19518 5788 19524 5840
rect 19576 5788 19582 5840
rect 8680 5732 9444 5760
rect 12176 5732 12756 5760
rect 4135 5666 4292 5694
rect 4341 5695 4399 5701
rect 4135 5663 4147 5666
rect 4089 5657 4147 5663
rect 4341 5661 4353 5695
rect 4387 5692 4399 5695
rect 6937 5695 6995 5701
rect 4387 5664 4752 5692
rect 4387 5661 4399 5664
rect 4341 5655 4399 5661
rect 4724 5636 4752 5664
rect 6937 5661 6949 5695
rect 6983 5692 6995 5695
rect 7116 5692 7144 5732
rect 6983 5664 7144 5692
rect 6983 5661 6995 5664
rect 6937 5655 6995 5661
rect 7190 5652 7196 5704
rect 7248 5652 7254 5704
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5692 7435 5695
rect 8386 5692 8392 5704
rect 7423 5664 8392 5692
rect 7423 5661 7435 5664
rect 7377 5655 7435 5661
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 8478 5652 8484 5704
rect 8536 5692 8542 5704
rect 8536 5664 9168 5692
rect 8536 5652 8542 5664
rect 1949 5627 2007 5633
rect 1596 5596 1900 5624
rect 1765 5559 1823 5565
rect 1765 5556 1777 5559
rect 1228 5528 1777 5556
rect 1765 5525 1777 5528
rect 1811 5525 1823 5559
rect 1872 5556 1900 5596
rect 1949 5593 1961 5627
rect 1995 5624 2007 5627
rect 3142 5624 3148 5636
rect 1995 5596 3148 5624
rect 1995 5593 2007 5596
rect 1949 5587 2007 5593
rect 3142 5584 3148 5596
rect 3200 5584 3206 5636
rect 3510 5584 3516 5636
rect 3568 5584 3574 5636
rect 4614 5633 4620 5636
rect 4586 5627 4620 5633
rect 4586 5593 4598 5627
rect 4586 5587 4620 5593
rect 4614 5584 4620 5587
rect 4672 5584 4678 5636
rect 4706 5584 4712 5636
rect 4764 5584 4770 5636
rect 6454 5624 6460 5636
rect 5736 5596 6460 5624
rect 2406 5556 2412 5568
rect 1872 5528 2412 5556
rect 1765 5519 1823 5525
rect 2406 5516 2412 5528
rect 2464 5516 2470 5568
rect 3053 5559 3111 5565
rect 3053 5525 3065 5559
rect 3099 5556 3111 5559
rect 3878 5556 3884 5568
rect 3099 5528 3884 5556
rect 3099 5525 3111 5528
rect 3053 5519 3111 5525
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 3970 5516 3976 5568
rect 4028 5556 4034 5568
rect 5074 5556 5080 5568
rect 4028 5528 5080 5556
rect 4028 5516 4034 5528
rect 5074 5516 5080 5528
rect 5132 5516 5138 5568
rect 5736 5565 5764 5596
rect 6454 5584 6460 5596
rect 6512 5584 6518 5636
rect 7622 5627 7680 5633
rect 7622 5624 7634 5627
rect 7392 5596 7634 5624
rect 7392 5568 7420 5596
rect 7622 5593 7634 5596
rect 7668 5593 7680 5627
rect 7622 5587 7680 5593
rect 5721 5559 5779 5565
rect 5721 5525 5733 5559
rect 5767 5525 5779 5559
rect 5721 5519 5779 5525
rect 5813 5559 5871 5565
rect 5813 5525 5825 5559
rect 5859 5556 5871 5559
rect 6822 5556 6828 5568
rect 5859 5528 6828 5556
rect 5859 5525 5871 5528
rect 5813 5519 5871 5525
rect 6822 5516 6828 5528
rect 6880 5516 6886 5568
rect 7374 5516 7380 5568
rect 7432 5516 7438 5568
rect 9140 5556 9168 5664
rect 9214 5652 9220 5704
rect 9272 5652 9278 5704
rect 9306 5652 9312 5704
rect 9364 5652 9370 5704
rect 9416 5692 9444 5732
rect 17678 5720 17684 5772
rect 17736 5760 17742 5772
rect 18693 5763 18751 5769
rect 18693 5760 18705 5763
rect 17736 5732 18705 5760
rect 17736 5720 17742 5732
rect 18693 5729 18705 5732
rect 18739 5729 18751 5763
rect 18693 5723 18751 5729
rect 19334 5720 19340 5772
rect 19392 5760 19398 5772
rect 20257 5763 20315 5769
rect 20257 5760 20269 5763
rect 19392 5732 20269 5760
rect 19392 5720 19398 5732
rect 20257 5729 20269 5732
rect 20303 5729 20315 5763
rect 20257 5723 20315 5729
rect 9416 5664 10364 5692
rect 9576 5627 9634 5633
rect 9576 5593 9588 5627
rect 9622 5593 9634 5627
rect 9576 5587 9634 5593
rect 9214 5556 9220 5568
rect 9140 5528 9220 5556
rect 9214 5516 9220 5528
rect 9272 5516 9278 5568
rect 9490 5516 9496 5568
rect 9548 5556 9554 5568
rect 9600 5556 9628 5587
rect 9548 5528 9628 5556
rect 10336 5556 10364 5664
rect 10778 5652 10784 5704
rect 10836 5652 10842 5704
rect 11054 5701 11060 5704
rect 11048 5692 11060 5701
rect 11015 5664 11060 5692
rect 11048 5655 11060 5664
rect 11054 5652 11060 5655
rect 11112 5652 11118 5704
rect 11330 5652 11336 5704
rect 11388 5692 11394 5704
rect 13725 5695 13783 5701
rect 11388 5664 12434 5692
rect 11388 5652 11394 5664
rect 10410 5584 10416 5636
rect 10468 5624 10474 5636
rect 12406 5624 12434 5664
rect 13725 5661 13737 5695
rect 13771 5692 13783 5695
rect 14182 5692 14188 5704
rect 13771 5664 14188 5692
rect 13771 5661 13783 5664
rect 13725 5655 13783 5661
rect 14182 5652 14188 5664
rect 14240 5652 14246 5704
rect 14829 5695 14887 5701
rect 14829 5661 14841 5695
rect 14875 5661 14887 5695
rect 14829 5655 14887 5661
rect 15013 5695 15071 5701
rect 15013 5661 15025 5695
rect 15059 5692 15071 5695
rect 15654 5692 15660 5704
rect 15059 5664 15660 5692
rect 15059 5661 15071 5664
rect 15013 5655 15071 5661
rect 13458 5627 13516 5633
rect 13458 5624 13470 5627
rect 10468 5596 12296 5624
rect 12406 5596 13470 5624
rect 10468 5584 10474 5596
rect 11698 5556 11704 5568
rect 10336 5528 11704 5556
rect 9548 5516 9554 5528
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 12268 5556 12296 5596
rect 13458 5593 13470 5596
rect 13504 5593 13516 5627
rect 13458 5587 13516 5593
rect 14553 5627 14611 5633
rect 14553 5593 14565 5627
rect 14599 5593 14611 5627
rect 14844 5624 14872 5655
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 16666 5652 16672 5704
rect 16724 5652 16730 5704
rect 18322 5692 18328 5704
rect 16868 5664 18328 5692
rect 15102 5624 15108 5636
rect 14844 5596 15108 5624
rect 14553 5587 14611 5593
rect 12345 5559 12403 5565
rect 12345 5556 12357 5559
rect 12268 5528 12357 5556
rect 12345 5525 12357 5528
rect 12391 5525 12403 5559
rect 14568 5556 14596 5587
rect 15102 5584 15108 5596
rect 15160 5584 15166 5636
rect 15280 5627 15338 5633
rect 15280 5593 15292 5627
rect 15326 5624 15338 5627
rect 15470 5624 15476 5636
rect 15326 5596 15476 5624
rect 15326 5593 15338 5596
rect 15280 5587 15338 5593
rect 15470 5584 15476 5596
rect 15528 5584 15534 5636
rect 15378 5556 15384 5568
rect 14568 5528 15384 5556
rect 12345 5519 12403 5525
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 16393 5559 16451 5565
rect 16393 5525 16405 5559
rect 16439 5556 16451 5559
rect 16868 5556 16896 5664
rect 18322 5652 18328 5664
rect 18380 5652 18386 5704
rect 19061 5695 19119 5701
rect 19061 5661 19073 5695
rect 19107 5661 19119 5695
rect 19061 5655 19119 5661
rect 16936 5627 16994 5633
rect 16936 5593 16948 5627
rect 16982 5624 16994 5627
rect 17402 5624 17408 5636
rect 16982 5596 17408 5624
rect 16982 5593 16994 5596
rect 16936 5587 16994 5593
rect 17402 5584 17408 5596
rect 17460 5584 17466 5636
rect 19076 5624 19104 5655
rect 19150 5652 19156 5704
rect 19208 5692 19214 5704
rect 19245 5695 19303 5701
rect 19245 5692 19257 5695
rect 19208 5664 19257 5692
rect 19208 5652 19214 5664
rect 19245 5661 19257 5664
rect 19291 5661 19303 5695
rect 19245 5655 19303 5661
rect 20162 5652 20168 5704
rect 20220 5652 20226 5704
rect 20364 5692 20392 5856
rect 20916 5769 20944 5856
rect 21008 5800 22876 5828
rect 20901 5763 20959 5769
rect 20901 5729 20913 5763
rect 20947 5729 20959 5763
rect 20901 5723 20959 5729
rect 21008 5692 21036 5800
rect 21450 5720 21456 5772
rect 21508 5760 21514 5772
rect 21545 5763 21603 5769
rect 21545 5760 21557 5763
rect 21508 5732 21557 5760
rect 21508 5720 21514 5732
rect 21545 5729 21557 5732
rect 21591 5729 21603 5763
rect 21545 5723 21603 5729
rect 21818 5720 21824 5772
rect 21876 5760 21882 5772
rect 21876 5732 22600 5760
rect 21876 5720 21882 5732
rect 22572 5701 22600 5732
rect 22848 5701 22876 5800
rect 20364 5664 21036 5692
rect 21913 5695 21971 5701
rect 21913 5661 21925 5695
rect 21959 5692 21971 5695
rect 22557 5695 22615 5701
rect 21959 5664 22508 5692
rect 21959 5661 21971 5664
rect 21913 5655 21971 5661
rect 21266 5624 21272 5636
rect 19076 5596 21272 5624
rect 21266 5584 21272 5596
rect 21324 5624 21330 5636
rect 21634 5624 21640 5636
rect 21324 5596 21640 5624
rect 21324 5584 21330 5596
rect 21634 5584 21640 5596
rect 21692 5584 21698 5636
rect 22480 5624 22508 5664
rect 22557 5661 22569 5695
rect 22603 5661 22615 5695
rect 22557 5655 22615 5661
rect 22833 5695 22891 5701
rect 22833 5661 22845 5695
rect 22879 5661 22891 5695
rect 22833 5655 22891 5661
rect 23290 5652 23296 5704
rect 23348 5652 23354 5704
rect 23382 5652 23388 5704
rect 23440 5652 23446 5704
rect 23400 5624 23428 5652
rect 22480 5596 23428 5624
rect 16439 5528 16896 5556
rect 16439 5525 16451 5528
rect 16393 5519 16451 5525
rect 18046 5516 18052 5568
rect 18104 5516 18110 5568
rect 1104 5466 23828 5488
rect 1104 5414 2658 5466
rect 2710 5414 2722 5466
rect 2774 5414 2786 5466
rect 2838 5414 2850 5466
rect 2902 5414 2914 5466
rect 2966 5414 2978 5466
rect 3030 5414 8658 5466
rect 8710 5414 8722 5466
rect 8774 5414 8786 5466
rect 8838 5414 8850 5466
rect 8902 5414 8914 5466
rect 8966 5414 8978 5466
rect 9030 5414 14658 5466
rect 14710 5414 14722 5466
rect 14774 5414 14786 5466
rect 14838 5414 14850 5466
rect 14902 5414 14914 5466
rect 14966 5414 14978 5466
rect 15030 5414 20658 5466
rect 20710 5414 20722 5466
rect 20774 5414 20786 5466
rect 20838 5414 20850 5466
rect 20902 5414 20914 5466
rect 20966 5414 20978 5466
rect 21030 5414 23828 5466
rect 1104 5392 23828 5414
rect 1946 5312 1952 5364
rect 2004 5312 2010 5364
rect 2041 5355 2099 5361
rect 2041 5321 2053 5355
rect 2087 5352 2099 5355
rect 2314 5352 2320 5364
rect 2087 5324 2320 5352
rect 2087 5321 2099 5324
rect 2041 5315 2099 5321
rect 2314 5312 2320 5324
rect 2372 5312 2378 5364
rect 3145 5355 3203 5361
rect 3145 5321 3157 5355
rect 3191 5352 3203 5355
rect 3694 5352 3700 5364
rect 3191 5324 3700 5352
rect 3191 5321 3203 5324
rect 3145 5315 3203 5321
rect 3694 5312 3700 5324
rect 3752 5312 3758 5364
rect 3786 5312 3792 5364
rect 3844 5312 3850 5364
rect 4614 5312 4620 5364
rect 4672 5352 4678 5364
rect 5721 5355 5779 5361
rect 5721 5352 5733 5355
rect 4672 5324 5733 5352
rect 4672 5312 4678 5324
rect 5721 5321 5733 5324
rect 5767 5321 5779 5355
rect 5721 5315 5779 5321
rect 6089 5355 6147 5361
rect 6089 5321 6101 5355
rect 6135 5352 6147 5355
rect 7282 5352 7288 5364
rect 6135 5324 7288 5352
rect 6135 5321 6147 5324
rect 6089 5315 6147 5321
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 9030 5312 9036 5364
rect 9088 5352 9094 5364
rect 9674 5352 9680 5364
rect 9088 5324 9680 5352
rect 9088 5312 9094 5324
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 10042 5312 10048 5364
rect 10100 5352 10106 5364
rect 13538 5352 13544 5364
rect 10100 5324 13544 5352
rect 10100 5312 10106 5324
rect 13538 5312 13544 5324
rect 13596 5312 13602 5364
rect 13814 5312 13820 5364
rect 13872 5312 13878 5364
rect 14182 5312 14188 5364
rect 14240 5352 14246 5364
rect 14645 5355 14703 5361
rect 14645 5352 14657 5355
rect 14240 5324 14657 5352
rect 14240 5312 14246 5324
rect 14645 5321 14657 5324
rect 14691 5321 14703 5355
rect 14645 5315 14703 5321
rect 15105 5355 15163 5361
rect 15105 5321 15117 5355
rect 15151 5352 15163 5355
rect 15286 5352 15292 5364
rect 15151 5324 15292 5352
rect 15151 5321 15163 5324
rect 15105 5315 15163 5321
rect 15286 5312 15292 5324
rect 15344 5312 15350 5364
rect 15654 5312 15660 5364
rect 15712 5312 15718 5364
rect 16022 5312 16028 5364
rect 16080 5352 16086 5364
rect 16301 5355 16359 5361
rect 16301 5352 16313 5355
rect 16080 5324 16313 5352
rect 16080 5312 16086 5324
rect 16301 5321 16313 5324
rect 16347 5321 16359 5355
rect 16301 5315 16359 5321
rect 17402 5312 17408 5364
rect 17460 5312 17466 5364
rect 18414 5312 18420 5364
rect 18472 5352 18478 5364
rect 18785 5355 18843 5361
rect 18785 5352 18797 5355
rect 18472 5324 18797 5352
rect 18472 5312 18478 5324
rect 18785 5321 18797 5324
rect 18831 5321 18843 5355
rect 18785 5315 18843 5321
rect 19150 5312 19156 5364
rect 19208 5312 19214 5364
rect 21266 5312 21272 5364
rect 21324 5312 21330 5364
rect 21358 5312 21364 5364
rect 21416 5312 21422 5364
rect 22189 5355 22247 5361
rect 22189 5321 22201 5355
rect 22235 5352 22247 5355
rect 22370 5352 22376 5364
rect 22235 5324 22376 5352
rect 22235 5321 22247 5324
rect 22189 5315 22247 5321
rect 22370 5312 22376 5324
rect 22428 5312 22434 5364
rect 23198 5312 23204 5364
rect 23256 5352 23262 5364
rect 23385 5355 23443 5361
rect 23385 5352 23397 5355
rect 23256 5324 23397 5352
rect 23256 5312 23262 5324
rect 23385 5321 23397 5324
rect 23431 5321 23443 5355
rect 23385 5315 23443 5321
rect 1964 5225 1992 5312
rect 3804 5284 3832 5312
rect 4157 5287 4215 5293
rect 3804 5256 4108 5284
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5216 3387 5219
rect 3970 5216 3976 5228
rect 3375 5188 3976 5216
rect 3375 5185 3387 5188
rect 3329 5179 3387 5185
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 4080 5225 4108 5256
rect 4157 5253 4169 5287
rect 4203 5284 4215 5287
rect 4203 5256 6408 5284
rect 4203 5253 4215 5256
rect 4157 5247 4215 5253
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 4430 5176 4436 5228
rect 4488 5216 4494 5228
rect 4597 5219 4655 5225
rect 4597 5216 4609 5219
rect 4488 5188 4609 5216
rect 4488 5176 4494 5188
rect 4597 5185 4609 5188
rect 4643 5185 4655 5219
rect 4597 5179 4655 5185
rect 4890 5176 4896 5228
rect 4948 5216 4954 5228
rect 5994 5216 6000 5228
rect 4948 5188 6000 5216
rect 4948 5176 4954 5188
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 6380 5225 6408 5256
rect 6454 5244 6460 5296
rect 6512 5284 6518 5296
rect 6610 5287 6668 5293
rect 6610 5284 6622 5287
rect 6512 5256 6622 5284
rect 6512 5244 6518 5256
rect 6610 5253 6622 5256
rect 6656 5253 6668 5287
rect 6610 5247 6668 5253
rect 8564 5287 8622 5293
rect 8564 5253 8576 5287
rect 8610 5284 8622 5287
rect 10410 5284 10416 5296
rect 8610 5256 10416 5284
rect 8610 5253 8622 5256
rect 8564 5247 8622 5253
rect 10410 5244 10416 5256
rect 10468 5244 10474 5296
rect 10502 5244 10508 5296
rect 10560 5284 10566 5296
rect 11066 5287 11124 5293
rect 11066 5284 11078 5287
rect 10560 5256 11078 5284
rect 10560 5244 10566 5256
rect 11066 5253 11078 5256
rect 11112 5253 11124 5287
rect 11066 5247 11124 5253
rect 12618 5244 12624 5296
rect 12676 5284 12682 5296
rect 13832 5284 13860 5312
rect 14921 5287 14979 5293
rect 14921 5284 14933 5287
rect 12676 5256 13584 5284
rect 13832 5256 14933 5284
rect 12676 5244 12682 5256
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 9398 5176 9404 5228
rect 9456 5216 9462 5228
rect 9766 5216 9772 5228
rect 9456 5188 9772 5216
rect 9456 5176 9462 5188
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 12894 5176 12900 5228
rect 12952 5216 12958 5228
rect 13458 5219 13516 5225
rect 13458 5216 13470 5219
rect 12952 5188 13470 5216
rect 12952 5176 12958 5188
rect 13458 5185 13470 5188
rect 13504 5185 13516 5219
rect 13556 5216 13584 5256
rect 14921 5253 14933 5256
rect 14967 5253 14979 5287
rect 19168 5284 19196 5312
rect 14921 5247 14979 5253
rect 16408 5256 19196 5284
rect 14369 5219 14427 5225
rect 14369 5216 14381 5219
rect 13556 5188 14381 5216
rect 13458 5179 13516 5185
rect 14369 5185 14381 5188
rect 14415 5185 14427 5219
rect 14369 5179 14427 5185
rect 14550 5176 14556 5228
rect 14608 5216 14614 5228
rect 14737 5219 14795 5225
rect 14737 5216 14749 5219
rect 14608 5188 14749 5216
rect 14608 5176 14614 5188
rect 14737 5185 14749 5188
rect 14783 5185 14795 5219
rect 14737 5179 14795 5185
rect 14829 5219 14887 5225
rect 14829 5185 14841 5219
rect 14875 5185 14887 5219
rect 14829 5179 14887 5185
rect 3510 5108 3516 5160
rect 3568 5148 3574 5160
rect 4341 5151 4399 5157
rect 4341 5148 4353 5151
rect 3568 5120 4353 5148
rect 3568 5108 3574 5120
rect 4341 5117 4353 5120
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 7374 5108 7380 5160
rect 7432 5148 7438 5160
rect 8297 5151 8355 5157
rect 8297 5148 8309 5151
rect 7432 5120 8309 5148
rect 7432 5108 7438 5120
rect 8297 5117 8309 5120
rect 8343 5117 8355 5151
rect 8297 5111 8355 5117
rect 11330 5108 11336 5160
rect 11388 5108 11394 5160
rect 13722 5108 13728 5160
rect 13780 5108 13786 5160
rect 14458 5108 14464 5160
rect 14516 5148 14522 5160
rect 14844 5148 14872 5179
rect 15194 5176 15200 5228
rect 15252 5216 15258 5228
rect 16408 5225 16436 5256
rect 15289 5219 15347 5225
rect 15289 5216 15301 5219
rect 15252 5188 15301 5216
rect 15252 5176 15258 5188
rect 15289 5185 15301 5188
rect 15335 5185 15347 5219
rect 15289 5179 15347 5185
rect 15749 5219 15807 5225
rect 15749 5185 15761 5219
rect 15795 5216 15807 5219
rect 16393 5219 16451 5225
rect 16393 5216 16405 5219
rect 15795 5188 16405 5216
rect 15795 5185 15807 5188
rect 15749 5179 15807 5185
rect 16393 5185 16405 5188
rect 16439 5185 16451 5219
rect 16393 5179 16451 5185
rect 16942 5176 16948 5228
rect 17000 5216 17006 5228
rect 17221 5219 17279 5225
rect 17221 5216 17233 5219
rect 17000 5188 17233 5216
rect 17000 5176 17006 5188
rect 17221 5185 17233 5188
rect 17267 5185 17279 5219
rect 17221 5179 17279 5185
rect 18141 5219 18199 5225
rect 18141 5185 18153 5219
rect 18187 5216 18199 5219
rect 18230 5216 18236 5228
rect 18187 5188 18236 5216
rect 18187 5185 18199 5188
rect 18141 5179 18199 5185
rect 18230 5176 18236 5188
rect 18288 5176 18294 5228
rect 18322 5176 18328 5228
rect 18380 5176 18386 5228
rect 18877 5219 18935 5225
rect 18877 5185 18889 5219
rect 18923 5216 18935 5219
rect 19058 5216 19064 5228
rect 18923 5188 19064 5216
rect 18923 5185 18935 5188
rect 18877 5179 18935 5185
rect 19058 5176 19064 5188
rect 19116 5176 19122 5228
rect 21284 5216 21312 5312
rect 21453 5219 21511 5225
rect 21453 5216 21465 5219
rect 21284 5188 21465 5216
rect 21453 5185 21465 5188
rect 21499 5185 21511 5219
rect 21453 5179 21511 5185
rect 22462 5176 22468 5228
rect 22520 5216 22526 5228
rect 22741 5219 22799 5225
rect 22741 5216 22753 5219
rect 22520 5188 22753 5216
rect 22520 5176 22526 5188
rect 22741 5185 22753 5188
rect 22787 5185 22799 5219
rect 22741 5179 22799 5185
rect 23293 5219 23351 5225
rect 23293 5185 23305 5219
rect 23339 5216 23351 5219
rect 23382 5216 23388 5228
rect 23339 5188 23388 5216
rect 23339 5185 23351 5188
rect 23293 5179 23351 5185
rect 23382 5176 23388 5188
rect 23440 5176 23446 5228
rect 14516 5120 14872 5148
rect 14516 5108 14522 5120
rect 15838 5108 15844 5160
rect 15896 5148 15902 5160
rect 16669 5151 16727 5157
rect 16669 5148 16681 5151
rect 15896 5120 16681 5148
rect 15896 5108 15902 5120
rect 16669 5117 16681 5120
rect 16715 5117 16727 5151
rect 16669 5111 16727 5117
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5148 18107 5151
rect 18340 5148 18368 5176
rect 18095 5120 18368 5148
rect 18095 5117 18107 5120
rect 18049 5111 18107 5117
rect 19426 5108 19432 5160
rect 19484 5108 19490 5160
rect 11698 5040 11704 5092
rect 11756 5080 11762 5092
rect 12345 5083 12403 5089
rect 12345 5080 12357 5083
rect 11756 5052 12357 5080
rect 11756 5040 11762 5052
rect 12345 5049 12357 5052
rect 12391 5049 12403 5083
rect 12345 5043 12403 5049
rect 18325 5083 18383 5089
rect 18325 5049 18337 5083
rect 18371 5080 18383 5083
rect 19444 5080 19472 5108
rect 18371 5052 19472 5080
rect 18371 5049 18383 5052
rect 18325 5043 18383 5049
rect 7742 4972 7748 5024
rect 7800 4972 7806 5024
rect 9674 4972 9680 5024
rect 9732 4972 9738 5024
rect 9953 5015 10011 5021
rect 9953 4981 9965 5015
rect 9999 5012 10011 5015
rect 10226 5012 10232 5024
rect 9999 4984 10232 5012
rect 9999 4981 10011 4984
rect 9953 4975 10011 4981
rect 10226 4972 10232 4984
rect 10284 5012 10290 5024
rect 10686 5012 10692 5024
rect 10284 4984 10692 5012
rect 10284 4972 10290 4984
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 12986 4972 12992 5024
rect 13044 5012 13050 5024
rect 13817 5015 13875 5021
rect 13817 5012 13829 5015
rect 13044 4984 13829 5012
rect 13044 4972 13050 4984
rect 13817 4981 13829 4984
rect 13863 4981 13875 5015
rect 13817 4975 13875 4981
rect 1104 4922 23828 4944
rect 1104 4870 1918 4922
rect 1970 4870 1982 4922
rect 2034 4870 2046 4922
rect 2098 4870 2110 4922
rect 2162 4870 2174 4922
rect 2226 4870 2238 4922
rect 2290 4870 7918 4922
rect 7970 4870 7982 4922
rect 8034 4870 8046 4922
rect 8098 4870 8110 4922
rect 8162 4870 8174 4922
rect 8226 4870 8238 4922
rect 8290 4870 13918 4922
rect 13970 4870 13982 4922
rect 14034 4870 14046 4922
rect 14098 4870 14110 4922
rect 14162 4870 14174 4922
rect 14226 4870 14238 4922
rect 14290 4870 19918 4922
rect 19970 4870 19982 4922
rect 20034 4870 20046 4922
rect 20098 4870 20110 4922
rect 20162 4870 20174 4922
rect 20226 4870 20238 4922
rect 20290 4870 23828 4922
rect 1104 4848 23828 4870
rect 5810 4768 5816 4820
rect 5868 4768 5874 4820
rect 6089 4811 6147 4817
rect 6089 4777 6101 4811
rect 6135 4808 6147 4811
rect 7374 4808 7380 4820
rect 6135 4780 7380 4808
rect 6135 4777 6147 4780
rect 6089 4771 6147 4777
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 7558 4768 7564 4820
rect 7616 4768 7622 4820
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 11241 4811 11299 4817
rect 11241 4808 11253 4811
rect 9640 4780 11253 4808
rect 9640 4768 9646 4780
rect 11241 4777 11253 4780
rect 11287 4777 11299 4811
rect 11241 4771 11299 4777
rect 13078 4768 13084 4820
rect 13136 4768 13142 4820
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 14277 4811 14335 4817
rect 14277 4808 14289 4811
rect 13872 4780 14289 4808
rect 13872 4768 13878 4780
rect 14277 4777 14289 4780
rect 14323 4777 14335 4811
rect 14277 4771 14335 4777
rect 16666 4768 16672 4820
rect 16724 4808 16730 4820
rect 16853 4811 16911 4817
rect 16853 4808 16865 4811
rect 16724 4780 16865 4808
rect 16724 4768 16730 4780
rect 16853 4777 16865 4780
rect 16899 4777 16911 4811
rect 16853 4771 16911 4777
rect 17126 4768 17132 4820
rect 17184 4768 17190 4820
rect 21726 4768 21732 4820
rect 21784 4768 21790 4820
rect 22738 4768 22744 4820
rect 22796 4808 22802 4820
rect 22833 4811 22891 4817
rect 22833 4808 22845 4811
rect 22796 4780 22845 4808
rect 22796 4768 22802 4780
rect 22833 4777 22845 4780
rect 22879 4777 22891 4811
rect 22833 4771 22891 4777
rect 6457 4743 6515 4749
rect 6457 4709 6469 4743
rect 6503 4740 6515 4743
rect 7576 4740 7604 4768
rect 6503 4712 7604 4740
rect 6503 4709 6515 4712
rect 6457 4703 6515 4709
rect 9398 4700 9404 4752
rect 9456 4700 9462 4752
rect 4062 4632 4068 4684
rect 4120 4672 4126 4684
rect 9493 4675 9551 4681
rect 4120 4644 9168 4672
rect 4120 4632 4126 4644
rect 5920 4613 5948 4644
rect 5905 4607 5963 4613
rect 5905 4573 5917 4607
rect 5951 4573 5963 4607
rect 5905 4567 5963 4573
rect 5994 4564 6000 4616
rect 6052 4564 6058 4616
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4604 6423 4607
rect 6411 4576 6592 4604
rect 6411 4573 6423 4576
rect 6365 4567 6423 4573
rect 6564 4536 6592 4576
rect 6638 4564 6644 4616
rect 6696 4564 6702 4616
rect 6730 4564 6736 4616
rect 6788 4564 6794 4616
rect 7098 4564 7104 4616
rect 7156 4604 7162 4616
rect 7285 4607 7343 4613
rect 7285 4604 7297 4607
rect 7156 4576 7297 4604
rect 7156 4564 7162 4576
rect 7285 4573 7297 4576
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4604 7435 4607
rect 7650 4604 7656 4616
rect 7423 4576 7656 4604
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 7650 4564 7656 4576
rect 7708 4564 7714 4616
rect 7742 4564 7748 4616
rect 7800 4604 7806 4616
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 7800 4576 7941 4604
rect 7800 4564 7806 4576
rect 7929 4573 7941 4576
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 8665 4607 8723 4613
rect 8665 4604 8677 4607
rect 8352 4576 8677 4604
rect 8352 4564 8358 4576
rect 8665 4573 8677 4576
rect 8711 4573 8723 4607
rect 8665 4567 8723 4573
rect 9030 4564 9036 4616
rect 9088 4564 9094 4616
rect 9140 4604 9168 4644
rect 9493 4641 9505 4675
rect 9539 4672 9551 4675
rect 9858 4672 9864 4684
rect 9539 4644 9864 4672
rect 9539 4641 9551 4644
rect 9493 4635 9551 4641
rect 9858 4632 9864 4644
rect 9916 4632 9922 4684
rect 9950 4632 9956 4684
rect 10008 4632 10014 4684
rect 12897 4675 12955 4681
rect 12897 4641 12909 4675
rect 12943 4672 12955 4675
rect 13357 4675 13415 4681
rect 13357 4672 13369 4675
rect 12943 4644 13369 4672
rect 12943 4641 12955 4644
rect 12897 4635 12955 4641
rect 13357 4641 13369 4644
rect 13403 4641 13415 4675
rect 17144 4672 17172 4768
rect 13357 4635 13415 4641
rect 14476 4644 17172 4672
rect 9968 4604 9996 4632
rect 10965 4607 11023 4613
rect 10965 4604 10977 4607
rect 9140 4576 9674 4604
rect 9968 4576 10977 4604
rect 6748 4536 6776 4564
rect 8478 4536 8484 4548
rect 6564 4508 8484 4536
rect 8478 4496 8484 4508
rect 8536 4496 8542 4548
rect 8110 4428 8116 4480
rect 8168 4428 8174 4480
rect 9048 4468 9076 4564
rect 9646 4536 9674 4576
rect 10965 4573 10977 4576
rect 11011 4573 11023 4607
rect 10965 4567 11023 4573
rect 11422 4564 11428 4616
rect 11480 4564 11486 4616
rect 12641 4607 12699 4613
rect 12641 4573 12653 4607
rect 12687 4604 12699 4607
rect 12986 4604 12992 4616
rect 12687 4576 12992 4604
rect 12687 4573 12699 4576
rect 12641 4567 12699 4573
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 13170 4564 13176 4616
rect 13228 4604 13234 4616
rect 13449 4607 13507 4613
rect 13228 4576 13400 4604
rect 13228 4564 13234 4576
rect 10042 4536 10048 4548
rect 9646 4508 10048 4536
rect 10042 4496 10048 4508
rect 10100 4496 10106 4548
rect 10318 4496 10324 4548
rect 10376 4536 10382 4548
rect 10698 4539 10756 4545
rect 10698 4536 10710 4539
rect 10376 4508 10710 4536
rect 10376 4496 10382 4508
rect 10698 4505 10710 4508
rect 10744 4505 10756 4539
rect 13372 4536 13400 4576
rect 13449 4573 13461 4607
rect 13495 4604 13507 4607
rect 13538 4604 13544 4616
rect 13495 4576 13544 4604
rect 13495 4573 13507 4576
rect 13449 4567 13507 4573
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 14476 4613 14504 4644
rect 22094 4632 22100 4684
rect 22152 4672 22158 4684
rect 22281 4675 22339 4681
rect 22281 4672 22293 4675
rect 22152 4644 22293 4672
rect 22152 4632 22158 4644
rect 22281 4641 22293 4644
rect 22327 4641 22339 4675
rect 22281 4635 22339 4641
rect 23474 4632 23480 4684
rect 23532 4632 23538 4684
rect 14461 4607 14519 4613
rect 14461 4573 14473 4607
rect 14507 4573 14519 4607
rect 14461 4567 14519 4573
rect 14550 4564 14556 4616
rect 14608 4564 14614 4616
rect 16945 4607 17003 4613
rect 16945 4573 16957 4607
rect 16991 4604 17003 4607
rect 19058 4604 19064 4616
rect 16991 4576 19064 4604
rect 16991 4573 17003 4576
rect 16945 4567 17003 4573
rect 19058 4564 19064 4576
rect 19116 4564 19122 4616
rect 14568 4536 14596 4564
rect 13372 4508 14596 4536
rect 10698 4499 10756 4505
rect 9490 4468 9496 4480
rect 9048 4440 9496 4468
rect 9490 4428 9496 4440
rect 9548 4428 9554 4480
rect 9582 4428 9588 4480
rect 9640 4428 9646 4480
rect 11517 4471 11575 4477
rect 11517 4437 11529 4471
rect 11563 4468 11575 4471
rect 12250 4468 12256 4480
rect 11563 4440 12256 4468
rect 11563 4437 11575 4440
rect 11517 4431 11575 4437
rect 12250 4428 12256 4440
rect 12308 4428 12314 4480
rect 1104 4378 23828 4400
rect 1104 4326 2658 4378
rect 2710 4326 2722 4378
rect 2774 4326 2786 4378
rect 2838 4326 2850 4378
rect 2902 4326 2914 4378
rect 2966 4326 2978 4378
rect 3030 4326 8658 4378
rect 8710 4326 8722 4378
rect 8774 4326 8786 4378
rect 8838 4326 8850 4378
rect 8902 4326 8914 4378
rect 8966 4326 8978 4378
rect 9030 4326 14658 4378
rect 14710 4326 14722 4378
rect 14774 4326 14786 4378
rect 14838 4326 14850 4378
rect 14902 4326 14914 4378
rect 14966 4326 14978 4378
rect 15030 4326 20658 4378
rect 20710 4326 20722 4378
rect 20774 4326 20786 4378
rect 20838 4326 20850 4378
rect 20902 4326 20914 4378
rect 20966 4326 20978 4378
rect 21030 4326 23828 4378
rect 1104 4304 23828 4326
rect 5994 4224 6000 4276
rect 6052 4224 6058 4276
rect 8110 4224 8116 4276
rect 8168 4224 8174 4276
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 9030 4264 9036 4276
rect 8352 4236 9036 4264
rect 8352 4224 8358 4236
rect 9030 4224 9036 4236
rect 9088 4224 9094 4276
rect 9585 4267 9643 4273
rect 9585 4233 9597 4267
rect 9631 4264 9643 4267
rect 9766 4264 9772 4276
rect 9631 4236 9772 4264
rect 9631 4233 9643 4236
rect 9585 4227 9643 4233
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 13081 4267 13139 4273
rect 13081 4233 13093 4267
rect 13127 4264 13139 4267
rect 13722 4264 13728 4276
rect 13127 4236 13728 4264
rect 13127 4233 13139 4236
rect 13081 4227 13139 4233
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 3418 4088 3424 4140
rect 3476 4088 3482 4140
rect 6012 4128 6040 4224
rect 6454 4128 6460 4140
rect 6012 4100 6460 4128
rect 6454 4088 6460 4100
rect 6512 4088 6518 4140
rect 6546 4088 6552 4140
rect 6604 4088 6610 4140
rect 6914 4088 6920 4140
rect 6972 4088 6978 4140
rect 7101 4131 7159 4137
rect 7101 4097 7113 4131
rect 7147 4128 7159 4131
rect 8128 4128 8156 4224
rect 12618 4156 12624 4208
rect 12676 4205 12682 4208
rect 12676 4196 12688 4205
rect 12676 4168 12721 4196
rect 12676 4159 12688 4168
rect 12676 4156 12682 4159
rect 13170 4156 13176 4208
rect 13228 4156 13234 4208
rect 7147 4100 8156 4128
rect 8389 4131 8447 4137
rect 7147 4097 7159 4100
rect 7101 4091 7159 4097
rect 8389 4097 8401 4131
rect 8435 4128 8447 4131
rect 8570 4128 8576 4140
rect 8435 4100 8576 4128
rect 8435 4097 8447 4100
rect 8389 4091 8447 4097
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 8849 4131 8907 4137
rect 8849 4097 8861 4131
rect 8895 4128 8907 4131
rect 9677 4131 9735 4137
rect 9677 4128 9689 4131
rect 8895 4100 9689 4128
rect 8895 4097 8907 4100
rect 8849 4091 8907 4097
rect 9677 4097 9689 4100
rect 9723 4097 9735 4131
rect 9677 4091 9735 4097
rect 9858 4088 9864 4140
rect 9916 4128 9922 4140
rect 10229 4131 10287 4137
rect 10229 4128 10241 4131
rect 9916 4100 10241 4128
rect 9916 4088 9922 4100
rect 10229 4097 10241 4100
rect 10275 4097 10287 4131
rect 10229 4091 10287 4097
rect 10413 4131 10471 4137
rect 10413 4097 10425 4131
rect 10459 4097 10471 4131
rect 10413 4091 10471 4097
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 10778 4128 10784 4140
rect 10551 4100 10784 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 3436 3992 3464 4088
rect 6932 4060 6960 4088
rect 7377 4063 7435 4069
rect 7377 4060 7389 4063
rect 6932 4032 7389 4060
rect 7377 4029 7389 4032
rect 7423 4029 7435 4063
rect 7377 4023 7435 4029
rect 9033 4063 9091 4069
rect 9033 4029 9045 4063
rect 9079 4060 9091 4063
rect 9214 4060 9220 4072
rect 9079 4032 9220 4060
rect 9079 4029 9091 4032
rect 9033 4023 9091 4029
rect 9214 4020 9220 4032
rect 9272 4020 9278 4072
rect 10428 4060 10456 4091
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 11238 4088 11244 4140
rect 11296 4128 11302 4140
rect 11333 4131 11391 4137
rect 11333 4128 11345 4131
rect 11296 4100 11345 4128
rect 11296 4088 11302 4100
rect 11333 4097 11345 4100
rect 11379 4097 11391 4131
rect 11333 4091 11391 4097
rect 11882 4088 11888 4140
rect 11940 4088 11946 4140
rect 13188 4127 13216 4156
rect 13173 4121 13231 4127
rect 10428 4032 10548 4060
rect 8297 3995 8355 4001
rect 8297 3992 8309 3995
rect 3436 3964 8309 3992
rect 8297 3961 8309 3964
rect 8343 3961 8355 3995
rect 10520 3992 10548 4032
rect 10686 4020 10692 4072
rect 10744 4020 10750 4072
rect 11054 3992 11060 4004
rect 10520 3964 11060 3992
rect 8297 3955 8355 3961
rect 11054 3952 11060 3964
rect 11112 3992 11118 4004
rect 11900 3992 11928 4088
rect 13173 4087 13185 4121
rect 13219 4087 13231 4121
rect 22554 4088 22560 4140
rect 22612 4088 22618 4140
rect 23106 4088 23112 4140
rect 23164 4128 23170 4140
rect 23201 4131 23259 4137
rect 23201 4128 23213 4131
rect 23164 4100 23213 4128
rect 23164 4088 23170 4100
rect 23201 4097 23213 4100
rect 23247 4097 23259 4131
rect 23201 4091 23259 4097
rect 13173 4081 13231 4087
rect 12897 4063 12955 4069
rect 12897 4029 12909 4063
rect 12943 4029 12955 4063
rect 12897 4023 12955 4029
rect 11112 3964 11928 3992
rect 12912 3992 12940 4023
rect 14366 3992 14372 4004
rect 12912 3964 14372 3992
rect 11112 3952 11118 3964
rect 14366 3952 14372 3964
rect 14424 3952 14430 4004
rect 7282 3884 7288 3936
rect 7340 3884 7346 3936
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3924 8079 3927
rect 8570 3924 8576 3936
rect 8067 3896 8576 3924
rect 8067 3893 8079 3896
rect 8021 3887 8079 3893
rect 8570 3884 8576 3896
rect 8628 3884 8634 3936
rect 8665 3927 8723 3933
rect 8665 3893 8677 3927
rect 8711 3924 8723 3927
rect 9122 3924 9128 3936
rect 8711 3896 9128 3924
rect 8711 3893 8723 3896
rect 8665 3887 8723 3893
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 11517 3927 11575 3933
rect 11517 3893 11529 3927
rect 11563 3924 11575 3927
rect 12894 3924 12900 3936
rect 11563 3896 12900 3924
rect 11563 3893 11575 3896
rect 11517 3887 11575 3893
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 1104 3834 23828 3856
rect 1104 3782 1918 3834
rect 1970 3782 1982 3834
rect 2034 3782 2046 3834
rect 2098 3782 2110 3834
rect 2162 3782 2174 3834
rect 2226 3782 2238 3834
rect 2290 3782 7918 3834
rect 7970 3782 7982 3834
rect 8034 3782 8046 3834
rect 8098 3782 8110 3834
rect 8162 3782 8174 3834
rect 8226 3782 8238 3834
rect 8290 3782 13918 3834
rect 13970 3782 13982 3834
rect 14034 3782 14046 3834
rect 14098 3782 14110 3834
rect 14162 3782 14174 3834
rect 14226 3782 14238 3834
rect 14290 3782 19918 3834
rect 19970 3782 19982 3834
rect 20034 3782 20046 3834
rect 20098 3782 20110 3834
rect 20162 3782 20174 3834
rect 20226 3782 20238 3834
rect 20290 3782 23828 3834
rect 1104 3760 23828 3782
rect 7190 3680 7196 3732
rect 7248 3720 7254 3732
rect 7561 3723 7619 3729
rect 7561 3720 7573 3723
rect 7248 3692 7573 3720
rect 7248 3680 7254 3692
rect 7561 3689 7573 3692
rect 7607 3689 7619 3723
rect 7561 3683 7619 3689
rect 8386 3680 8392 3732
rect 8444 3720 8450 3732
rect 8665 3723 8723 3729
rect 8665 3720 8677 3723
rect 8444 3692 8677 3720
rect 8444 3680 8450 3692
rect 8665 3689 8677 3692
rect 8711 3689 8723 3723
rect 8665 3683 8723 3689
rect 9030 3680 9036 3732
rect 9088 3680 9094 3732
rect 9306 3680 9312 3732
rect 9364 3720 9370 3732
rect 10413 3723 10471 3729
rect 10413 3720 10425 3723
rect 9364 3692 10425 3720
rect 9364 3680 9370 3692
rect 10413 3689 10425 3692
rect 10459 3689 10471 3723
rect 10413 3683 10471 3689
rect 11330 3680 11336 3732
rect 11388 3720 11394 3732
rect 11885 3723 11943 3729
rect 11885 3720 11897 3723
rect 11388 3692 11897 3720
rect 11388 3680 11394 3692
rect 11885 3689 11897 3692
rect 11931 3689 11943 3723
rect 11885 3683 11943 3689
rect 12434 3680 12440 3732
rect 12492 3680 12498 3732
rect 7466 3612 7472 3664
rect 7524 3612 7530 3664
rect 8570 3612 8576 3664
rect 8628 3652 8634 3664
rect 9125 3655 9183 3661
rect 9125 3652 9137 3655
rect 8628 3624 9137 3652
rect 8628 3612 8634 3624
rect 9125 3621 9137 3624
rect 9171 3621 9183 3655
rect 9125 3615 9183 3621
rect 9398 3612 9404 3664
rect 9456 3652 9462 3664
rect 9585 3655 9643 3661
rect 9585 3652 9597 3655
rect 9456 3624 9597 3652
rect 9456 3612 9462 3624
rect 9585 3621 9597 3624
rect 9631 3621 9643 3655
rect 9585 3615 9643 3621
rect 11514 3612 11520 3664
rect 11572 3612 11578 3664
rect 7484 3584 7512 3612
rect 12161 3587 12219 3593
rect 12161 3584 12173 3587
rect 7484 3556 12173 3584
rect 12161 3553 12173 3556
rect 12207 3553 12219 3587
rect 12161 3547 12219 3553
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 7653 3519 7711 3525
rect 7653 3516 7665 3519
rect 6512 3488 7665 3516
rect 6512 3476 6518 3488
rect 7653 3485 7665 3488
rect 7699 3485 7711 3519
rect 7653 3479 7711 3485
rect 7668 3448 7696 3479
rect 8478 3476 8484 3528
rect 8536 3516 8542 3528
rect 8757 3519 8815 3525
rect 8757 3516 8769 3519
rect 8536 3488 8769 3516
rect 8536 3476 8542 3488
rect 8757 3485 8769 3488
rect 8803 3485 8815 3519
rect 8757 3479 8815 3485
rect 9490 3476 9496 3528
rect 9548 3476 9554 3528
rect 9674 3476 9680 3528
rect 9732 3516 9738 3528
rect 10137 3519 10195 3525
rect 10137 3516 10149 3519
rect 9732 3488 10149 3516
rect 9732 3476 9738 3488
rect 10137 3485 10149 3488
rect 10183 3485 10195 3519
rect 10137 3479 10195 3485
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3516 10563 3519
rect 11054 3516 11060 3528
rect 10551 3488 11060 3516
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 11606 3476 11612 3528
rect 11664 3516 11670 3528
rect 11701 3519 11759 3525
rect 11701 3516 11713 3519
rect 11664 3488 11713 3516
rect 11664 3476 11670 3488
rect 11701 3485 11713 3488
rect 11747 3485 11759 3519
rect 11701 3479 11759 3485
rect 11974 3476 11980 3528
rect 12032 3476 12038 3528
rect 12069 3519 12127 3525
rect 12069 3485 12081 3519
rect 12115 3485 12127 3519
rect 12069 3479 12127 3485
rect 12529 3519 12587 3525
rect 12529 3485 12541 3519
rect 12575 3516 12587 3519
rect 13538 3516 13544 3528
rect 12575 3488 13544 3516
rect 12575 3485 12587 3488
rect 12529 3479 12587 3485
rect 12084 3448 12112 3479
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 7668 3420 12112 3448
rect 1104 3290 23828 3312
rect 1104 3238 2658 3290
rect 2710 3238 2722 3290
rect 2774 3238 2786 3290
rect 2838 3238 2850 3290
rect 2902 3238 2914 3290
rect 2966 3238 2978 3290
rect 3030 3238 8658 3290
rect 8710 3238 8722 3290
rect 8774 3238 8786 3290
rect 8838 3238 8850 3290
rect 8902 3238 8914 3290
rect 8966 3238 8978 3290
rect 9030 3238 14658 3290
rect 14710 3238 14722 3290
rect 14774 3238 14786 3290
rect 14838 3238 14850 3290
rect 14902 3238 14914 3290
rect 14966 3238 14978 3290
rect 15030 3238 20658 3290
rect 20710 3238 20722 3290
rect 20774 3238 20786 3290
rect 20838 3238 20850 3290
rect 20902 3238 20914 3290
rect 20966 3238 20978 3290
rect 21030 3238 23828 3290
rect 1104 3216 23828 3238
rect 6362 3000 6368 3052
rect 6420 3040 6426 3052
rect 11609 3043 11667 3049
rect 11609 3040 11621 3043
rect 6420 3012 11621 3040
rect 6420 3000 6426 3012
rect 11609 3009 11621 3012
rect 11655 3009 11667 3043
rect 11609 3003 11667 3009
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 11885 2975 11943 2981
rect 11885 2972 11897 2975
rect 11020 2944 11897 2972
rect 11020 2932 11026 2944
rect 11885 2941 11897 2944
rect 11931 2941 11943 2975
rect 11885 2935 11943 2941
rect 1104 2746 23828 2768
rect 1104 2694 1918 2746
rect 1970 2694 1982 2746
rect 2034 2694 2046 2746
rect 2098 2694 2110 2746
rect 2162 2694 2174 2746
rect 2226 2694 2238 2746
rect 2290 2694 7918 2746
rect 7970 2694 7982 2746
rect 8034 2694 8046 2746
rect 8098 2694 8110 2746
rect 8162 2694 8174 2746
rect 8226 2694 8238 2746
rect 8290 2694 13918 2746
rect 13970 2694 13982 2746
rect 14034 2694 14046 2746
rect 14098 2694 14110 2746
rect 14162 2694 14174 2746
rect 14226 2694 14238 2746
rect 14290 2694 19918 2746
rect 19970 2694 19982 2746
rect 20034 2694 20046 2746
rect 20098 2694 20110 2746
rect 20162 2694 20174 2746
rect 20226 2694 20238 2746
rect 20290 2694 23828 2746
rect 1104 2672 23828 2694
rect 6270 2524 6276 2576
rect 6328 2564 6334 2576
rect 6328 2536 7972 2564
rect 6328 2524 6334 2536
rect 7190 2456 7196 2508
rect 7248 2496 7254 2508
rect 7377 2499 7435 2505
rect 7377 2496 7389 2499
rect 7248 2468 7389 2496
rect 7248 2456 7254 2468
rect 7377 2465 7389 2468
rect 7423 2465 7435 2499
rect 7377 2459 7435 2465
rect 5442 2388 5448 2440
rect 5500 2428 5506 2440
rect 7944 2437 7972 2536
rect 10689 2499 10747 2505
rect 10689 2465 10701 2499
rect 10735 2496 10747 2499
rect 11790 2496 11796 2508
rect 10735 2468 11796 2496
rect 10735 2465 10747 2468
rect 10689 2459 10747 2465
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 12268 2468 13032 2496
rect 12268 2440 12296 2468
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 5500 2400 7113 2428
rect 5500 2388 5506 2400
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 10410 2388 10416 2440
rect 10468 2388 10474 2440
rect 12250 2388 12256 2440
rect 12308 2388 12314 2440
rect 12526 2388 12532 2440
rect 12584 2388 12590 2440
rect 13004 2437 13032 2468
rect 12989 2431 13047 2437
rect 12989 2397 13001 2431
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 13354 2388 13360 2440
rect 13412 2428 13418 2440
rect 14185 2431 14243 2437
rect 14185 2428 14197 2431
rect 13412 2400 14197 2428
rect 13412 2388 13418 2400
rect 14185 2397 14197 2400
rect 14231 2397 14243 2431
rect 14185 2391 14243 2397
rect 17034 2388 17040 2440
rect 17092 2428 17098 2440
rect 17681 2431 17739 2437
rect 17681 2428 17693 2431
rect 17092 2400 17693 2428
rect 17092 2388 17098 2400
rect 17681 2397 17693 2400
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 18230 2388 18236 2440
rect 18288 2388 18294 2440
rect 7742 2320 7748 2372
rect 7800 2360 7806 2372
rect 8297 2363 8355 2369
rect 8297 2360 8309 2363
rect 7800 2332 8309 2360
rect 7800 2320 7806 2332
rect 8297 2329 8309 2332
rect 8343 2329 8355 2363
rect 8297 2323 8355 2329
rect 12158 2320 12164 2372
rect 12216 2320 12222 2372
rect 12894 2320 12900 2372
rect 12952 2360 12958 2372
rect 13265 2363 13323 2369
rect 13265 2360 13277 2363
rect 12952 2332 13277 2360
rect 12952 2320 12958 2332
rect 13265 2329 13277 2332
rect 13311 2329 13323 2363
rect 13265 2323 13323 2329
rect 13538 2320 13544 2372
rect 13596 2360 13602 2372
rect 14553 2363 14611 2369
rect 14553 2360 14565 2363
rect 13596 2332 14565 2360
rect 13596 2320 13602 2332
rect 14553 2329 14565 2332
rect 14599 2329 14611 2363
rect 14553 2323 14611 2329
rect 17310 2320 17316 2372
rect 17368 2320 17374 2372
rect 18046 2320 18052 2372
rect 18104 2360 18110 2372
rect 18601 2363 18659 2369
rect 18601 2360 18613 2363
rect 18104 2332 18613 2360
rect 18104 2320 18110 2332
rect 18601 2329 18613 2332
rect 18647 2329 18659 2363
rect 18601 2323 18659 2329
rect 1104 2202 23828 2224
rect 1104 2150 2658 2202
rect 2710 2150 2722 2202
rect 2774 2150 2786 2202
rect 2838 2150 2850 2202
rect 2902 2150 2914 2202
rect 2966 2150 2978 2202
rect 3030 2150 8658 2202
rect 8710 2150 8722 2202
rect 8774 2150 8786 2202
rect 8838 2150 8850 2202
rect 8902 2150 8914 2202
rect 8966 2150 8978 2202
rect 9030 2150 14658 2202
rect 14710 2150 14722 2202
rect 14774 2150 14786 2202
rect 14838 2150 14850 2202
rect 14902 2150 14914 2202
rect 14966 2150 14978 2202
rect 15030 2150 20658 2202
rect 20710 2150 20722 2202
rect 20774 2150 20786 2202
rect 20838 2150 20850 2202
rect 20902 2150 20914 2202
rect 20966 2150 20978 2202
rect 21030 2150 23828 2202
rect 1104 2128 23828 2150
<< via1 >>
rect 1918 24454 1970 24506
rect 1982 24454 2034 24506
rect 2046 24454 2098 24506
rect 2110 24454 2162 24506
rect 2174 24454 2226 24506
rect 2238 24454 2290 24506
rect 7918 24454 7970 24506
rect 7982 24454 8034 24506
rect 8046 24454 8098 24506
rect 8110 24454 8162 24506
rect 8174 24454 8226 24506
rect 8238 24454 8290 24506
rect 13918 24454 13970 24506
rect 13982 24454 14034 24506
rect 14046 24454 14098 24506
rect 14110 24454 14162 24506
rect 14174 24454 14226 24506
rect 14238 24454 14290 24506
rect 19918 24454 19970 24506
rect 19982 24454 20034 24506
rect 20046 24454 20098 24506
rect 20110 24454 20162 24506
rect 20174 24454 20226 24506
rect 20238 24454 20290 24506
rect 7748 24216 7800 24268
rect 8392 24216 8444 24268
rect 10968 24216 11020 24268
rect 13544 24216 13596 24268
rect 14464 24216 14516 24268
rect 7564 24148 7616 24200
rect 9588 24148 9640 24200
rect 10784 24148 10836 24200
rect 12992 24148 13044 24200
rect 14556 24148 14608 24200
rect 14832 24216 14884 24268
rect 15384 24148 15436 24200
rect 2658 23910 2710 23962
rect 2722 23910 2774 23962
rect 2786 23910 2838 23962
rect 2850 23910 2902 23962
rect 2914 23910 2966 23962
rect 2978 23910 3030 23962
rect 8658 23910 8710 23962
rect 8722 23910 8774 23962
rect 8786 23910 8838 23962
rect 8850 23910 8902 23962
rect 8914 23910 8966 23962
rect 8978 23910 9030 23962
rect 14658 23910 14710 23962
rect 14722 23910 14774 23962
rect 14786 23910 14838 23962
rect 14850 23910 14902 23962
rect 14914 23910 14966 23962
rect 14978 23910 15030 23962
rect 20658 23910 20710 23962
rect 20722 23910 20774 23962
rect 20786 23910 20838 23962
rect 20850 23910 20902 23962
rect 20914 23910 20966 23962
rect 20978 23910 21030 23962
rect 1918 23366 1970 23418
rect 1982 23366 2034 23418
rect 2046 23366 2098 23418
rect 2110 23366 2162 23418
rect 2174 23366 2226 23418
rect 2238 23366 2290 23418
rect 7918 23366 7970 23418
rect 7982 23366 8034 23418
rect 8046 23366 8098 23418
rect 8110 23366 8162 23418
rect 8174 23366 8226 23418
rect 8238 23366 8290 23418
rect 13918 23366 13970 23418
rect 13982 23366 14034 23418
rect 14046 23366 14098 23418
rect 14110 23366 14162 23418
rect 14174 23366 14226 23418
rect 14238 23366 14290 23418
rect 19918 23366 19970 23418
rect 19982 23366 20034 23418
rect 20046 23366 20098 23418
rect 20110 23366 20162 23418
rect 20174 23366 20226 23418
rect 20238 23366 20290 23418
rect 2658 22822 2710 22874
rect 2722 22822 2774 22874
rect 2786 22822 2838 22874
rect 2850 22822 2902 22874
rect 2914 22822 2966 22874
rect 2978 22822 3030 22874
rect 8658 22822 8710 22874
rect 8722 22822 8774 22874
rect 8786 22822 8838 22874
rect 8850 22822 8902 22874
rect 8914 22822 8966 22874
rect 8978 22822 9030 22874
rect 14658 22822 14710 22874
rect 14722 22822 14774 22874
rect 14786 22822 14838 22874
rect 14850 22822 14902 22874
rect 14914 22822 14966 22874
rect 14978 22822 15030 22874
rect 20658 22822 20710 22874
rect 20722 22822 20774 22874
rect 20786 22822 20838 22874
rect 20850 22822 20902 22874
rect 20914 22822 20966 22874
rect 20978 22822 21030 22874
rect 16488 22584 16540 22636
rect 10968 22380 11020 22432
rect 1918 22278 1970 22330
rect 1982 22278 2034 22330
rect 2046 22278 2098 22330
rect 2110 22278 2162 22330
rect 2174 22278 2226 22330
rect 2238 22278 2290 22330
rect 7918 22278 7970 22330
rect 7982 22278 8034 22330
rect 8046 22278 8098 22330
rect 8110 22278 8162 22330
rect 8174 22278 8226 22330
rect 8238 22278 8290 22330
rect 13918 22278 13970 22330
rect 13982 22278 14034 22330
rect 14046 22278 14098 22330
rect 14110 22278 14162 22330
rect 14174 22278 14226 22330
rect 14238 22278 14290 22330
rect 19918 22278 19970 22330
rect 19982 22278 20034 22330
rect 20046 22278 20098 22330
rect 20110 22278 20162 22330
rect 20174 22278 20226 22330
rect 20238 22278 20290 22330
rect 10324 22108 10376 22160
rect 10048 22040 10100 22092
rect 7840 21904 7892 21956
rect 6828 21836 6880 21888
rect 8576 21836 8628 21888
rect 9956 21972 10008 22024
rect 10508 21904 10560 21956
rect 10600 21904 10652 21956
rect 10968 21947 11020 21956
rect 10968 21913 11002 21947
rect 11002 21913 11020 21947
rect 10968 21904 11020 21913
rect 12624 22015 12676 22024
rect 12624 21981 12633 22015
rect 12633 21981 12667 22015
rect 12667 21981 12676 22015
rect 12624 21972 12676 21981
rect 14280 22015 14332 22024
rect 14280 21981 14289 22015
rect 14289 21981 14323 22015
rect 14323 21981 14332 22015
rect 14280 21972 14332 21981
rect 11060 21836 11112 21888
rect 12072 21879 12124 21888
rect 12072 21845 12081 21879
rect 12081 21845 12115 21879
rect 12115 21845 12124 21879
rect 12072 21836 12124 21845
rect 13176 21904 13228 21956
rect 13268 21879 13320 21888
rect 13268 21845 13277 21879
rect 13277 21845 13311 21879
rect 13311 21845 13320 21879
rect 13268 21836 13320 21845
rect 13728 21836 13780 21888
rect 13820 21836 13872 21888
rect 14464 21879 14516 21888
rect 14464 21845 14473 21879
rect 14473 21845 14507 21879
rect 14507 21845 14516 21879
rect 14464 21836 14516 21845
rect 15292 21879 15344 21888
rect 15292 21845 15301 21879
rect 15301 21845 15335 21879
rect 15335 21845 15344 21879
rect 15292 21836 15344 21845
rect 15476 21836 15528 21888
rect 2658 21734 2710 21786
rect 2722 21734 2774 21786
rect 2786 21734 2838 21786
rect 2850 21734 2902 21786
rect 2914 21734 2966 21786
rect 2978 21734 3030 21786
rect 8658 21734 8710 21786
rect 8722 21734 8774 21786
rect 8786 21734 8838 21786
rect 8850 21734 8902 21786
rect 8914 21734 8966 21786
rect 8978 21734 9030 21786
rect 14658 21734 14710 21786
rect 14722 21734 14774 21786
rect 14786 21734 14838 21786
rect 14850 21734 14902 21786
rect 14914 21734 14966 21786
rect 14978 21734 15030 21786
rect 20658 21734 20710 21786
rect 20722 21734 20774 21786
rect 20786 21734 20838 21786
rect 20850 21734 20902 21786
rect 20914 21734 20966 21786
rect 20978 21734 21030 21786
rect 10324 21675 10376 21684
rect 10324 21641 10333 21675
rect 10333 21641 10367 21675
rect 10367 21641 10376 21675
rect 10324 21632 10376 21641
rect 10508 21632 10560 21684
rect 11888 21632 11940 21684
rect 11060 21564 11112 21616
rect 13728 21564 13780 21616
rect 5632 21496 5684 21548
rect 10508 21496 10560 21548
rect 6552 21471 6604 21480
rect 6552 21437 6561 21471
rect 6561 21437 6595 21471
rect 6595 21437 6604 21471
rect 6552 21428 6604 21437
rect 7656 21428 7708 21480
rect 9496 21428 9548 21480
rect 9772 21471 9824 21480
rect 9772 21437 9781 21471
rect 9781 21437 9815 21471
rect 9815 21437 9824 21471
rect 9772 21428 9824 21437
rect 10416 21471 10468 21480
rect 10416 21437 10425 21471
rect 10425 21437 10459 21471
rect 10459 21437 10468 21471
rect 10416 21428 10468 21437
rect 11612 21496 11664 21548
rect 12624 21496 12676 21548
rect 15476 21539 15528 21548
rect 15476 21505 15485 21539
rect 15485 21505 15519 21539
rect 15519 21505 15528 21539
rect 15476 21496 15528 21505
rect 11796 21471 11848 21480
rect 11796 21437 11805 21471
rect 11805 21437 11839 21471
rect 11839 21437 11848 21471
rect 11796 21428 11848 21437
rect 14556 21471 14608 21480
rect 14556 21437 14565 21471
rect 14565 21437 14599 21471
rect 14599 21437 14608 21471
rect 14556 21428 14608 21437
rect 15568 21428 15620 21480
rect 17224 21471 17276 21480
rect 17224 21437 17233 21471
rect 17233 21437 17267 21471
rect 17267 21437 17276 21471
rect 17224 21428 17276 21437
rect 18144 21471 18196 21480
rect 18144 21437 18153 21471
rect 18153 21437 18187 21471
rect 18187 21437 18196 21471
rect 18144 21428 18196 21437
rect 7748 21292 7800 21344
rect 8484 21292 8536 21344
rect 9312 21292 9364 21344
rect 9404 21292 9456 21344
rect 11152 21292 11204 21344
rect 11244 21335 11296 21344
rect 11244 21301 11253 21335
rect 11253 21301 11287 21335
rect 11287 21301 11296 21335
rect 11244 21292 11296 21301
rect 11612 21335 11664 21344
rect 11612 21301 11621 21335
rect 11621 21301 11655 21335
rect 11655 21301 11664 21335
rect 11612 21292 11664 21301
rect 12440 21335 12492 21344
rect 12440 21301 12449 21335
rect 12449 21301 12483 21335
rect 12483 21301 12492 21335
rect 12440 21292 12492 21301
rect 13728 21292 13780 21344
rect 14740 21292 14792 21344
rect 15200 21335 15252 21344
rect 15200 21301 15209 21335
rect 15209 21301 15243 21335
rect 15243 21301 15252 21335
rect 15200 21292 15252 21301
rect 15384 21335 15436 21344
rect 15384 21301 15393 21335
rect 15393 21301 15427 21335
rect 15427 21301 15436 21335
rect 15384 21292 15436 21301
rect 16304 21335 16356 21344
rect 16304 21301 16313 21335
rect 16313 21301 16347 21335
rect 16347 21301 16356 21335
rect 16304 21292 16356 21301
rect 16672 21335 16724 21344
rect 16672 21301 16681 21335
rect 16681 21301 16715 21335
rect 16715 21301 16724 21335
rect 16672 21292 16724 21301
rect 18788 21335 18840 21344
rect 18788 21301 18797 21335
rect 18797 21301 18831 21335
rect 18831 21301 18840 21335
rect 18788 21292 18840 21301
rect 1918 21190 1970 21242
rect 1982 21190 2034 21242
rect 2046 21190 2098 21242
rect 2110 21190 2162 21242
rect 2174 21190 2226 21242
rect 2238 21190 2290 21242
rect 7918 21190 7970 21242
rect 7982 21190 8034 21242
rect 8046 21190 8098 21242
rect 8110 21190 8162 21242
rect 8174 21190 8226 21242
rect 8238 21190 8290 21242
rect 13918 21190 13970 21242
rect 13982 21190 14034 21242
rect 14046 21190 14098 21242
rect 14110 21190 14162 21242
rect 14174 21190 14226 21242
rect 14238 21190 14290 21242
rect 19918 21190 19970 21242
rect 19982 21190 20034 21242
rect 20046 21190 20098 21242
rect 20110 21190 20162 21242
rect 20174 21190 20226 21242
rect 20238 21190 20290 21242
rect 10968 21131 11020 21140
rect 10968 21097 10977 21131
rect 10977 21097 11011 21131
rect 11011 21097 11020 21131
rect 10968 21088 11020 21097
rect 5540 20952 5592 21004
rect 6184 20952 6236 21004
rect 6552 20952 6604 21004
rect 11244 21088 11296 21140
rect 12440 21088 12492 21140
rect 6736 20884 6788 20936
rect 4896 20816 4948 20868
rect 7840 20884 7892 20936
rect 14740 21088 14792 21140
rect 15292 21088 15344 21140
rect 15568 21088 15620 21140
rect 9220 20816 9272 20868
rect 10600 20816 10652 20868
rect 12532 20927 12584 20936
rect 12532 20893 12541 20927
rect 12541 20893 12575 20927
rect 12575 20893 12584 20927
rect 12532 20884 12584 20893
rect 13728 20884 13780 20936
rect 14648 20884 14700 20936
rect 16304 20884 16356 20936
rect 17776 20884 17828 20936
rect 18420 20884 18472 20936
rect 11336 20859 11388 20868
rect 11336 20825 11370 20859
rect 11370 20825 11388 20859
rect 11336 20816 11388 20825
rect 4344 20748 4396 20800
rect 5356 20748 5408 20800
rect 6920 20748 6972 20800
rect 7012 20748 7064 20800
rect 7840 20748 7892 20800
rect 8300 20748 8352 20800
rect 8392 20791 8444 20800
rect 8392 20757 8401 20791
rect 8401 20757 8435 20791
rect 8435 20757 8444 20791
rect 8392 20748 8444 20757
rect 9128 20748 9180 20800
rect 9404 20748 9456 20800
rect 11060 20748 11112 20800
rect 11796 20748 11848 20800
rect 19524 20816 19576 20868
rect 15568 20748 15620 20800
rect 18052 20791 18104 20800
rect 18052 20757 18061 20791
rect 18061 20757 18095 20791
rect 18095 20757 18104 20791
rect 18052 20748 18104 20757
rect 19340 20791 19392 20800
rect 19340 20757 19349 20791
rect 19349 20757 19383 20791
rect 19383 20757 19392 20791
rect 19340 20748 19392 20757
rect 2658 20646 2710 20698
rect 2722 20646 2774 20698
rect 2786 20646 2838 20698
rect 2850 20646 2902 20698
rect 2914 20646 2966 20698
rect 2978 20646 3030 20698
rect 8658 20646 8710 20698
rect 8722 20646 8774 20698
rect 8786 20646 8838 20698
rect 8850 20646 8902 20698
rect 8914 20646 8966 20698
rect 8978 20646 9030 20698
rect 14658 20646 14710 20698
rect 14722 20646 14774 20698
rect 14786 20646 14838 20698
rect 14850 20646 14902 20698
rect 14914 20646 14966 20698
rect 14978 20646 15030 20698
rect 20658 20646 20710 20698
rect 20722 20646 20774 20698
rect 20786 20646 20838 20698
rect 20850 20646 20902 20698
rect 20914 20646 20966 20698
rect 20978 20646 21030 20698
rect 4804 20451 4856 20460
rect 4804 20417 4813 20451
rect 4813 20417 4847 20451
rect 4847 20417 4856 20451
rect 4804 20408 4856 20417
rect 5356 20408 5408 20460
rect 5448 20408 5500 20460
rect 6644 20408 6696 20460
rect 8300 20544 8352 20596
rect 8668 20544 8720 20596
rect 10416 20544 10468 20596
rect 11336 20587 11388 20596
rect 11336 20553 11345 20587
rect 11345 20553 11379 20587
rect 11379 20553 11388 20587
rect 11336 20544 11388 20553
rect 7748 20408 7800 20460
rect 9312 20476 9364 20528
rect 11796 20519 11848 20528
rect 11796 20485 11830 20519
rect 11830 20485 11848 20519
rect 11796 20476 11848 20485
rect 8576 20408 8628 20460
rect 9588 20408 9640 20460
rect 14464 20544 14516 20596
rect 17224 20544 17276 20596
rect 9956 20383 10008 20392
rect 9956 20349 9965 20383
rect 9965 20349 9999 20383
rect 9999 20349 10008 20383
rect 9956 20340 10008 20349
rect 11520 20383 11572 20392
rect 11520 20349 11529 20383
rect 11529 20349 11563 20383
rect 11563 20349 11572 20383
rect 11520 20340 11572 20349
rect 15292 20476 15344 20528
rect 18144 20476 18196 20528
rect 18788 20476 18840 20528
rect 15200 20408 15252 20460
rect 18052 20408 18104 20460
rect 6276 20272 6328 20324
rect 14464 20272 14516 20324
rect 6368 20204 6420 20256
rect 6552 20247 6604 20256
rect 6552 20213 6561 20247
rect 6561 20213 6595 20247
rect 6595 20213 6604 20247
rect 6552 20204 6604 20213
rect 7656 20204 7708 20256
rect 15108 20204 15160 20256
rect 16672 20340 16724 20392
rect 17224 20383 17276 20392
rect 17224 20349 17233 20383
rect 17233 20349 17267 20383
rect 17267 20349 17276 20383
rect 17224 20340 17276 20349
rect 17408 20383 17460 20392
rect 17408 20349 17417 20383
rect 17417 20349 17451 20383
rect 17451 20349 17460 20383
rect 17408 20340 17460 20349
rect 16488 20247 16540 20256
rect 16488 20213 16497 20247
rect 16497 20213 16531 20247
rect 16531 20213 16540 20247
rect 16488 20204 16540 20213
rect 16672 20247 16724 20256
rect 16672 20213 16681 20247
rect 16681 20213 16715 20247
rect 16715 20213 16724 20247
rect 16672 20204 16724 20213
rect 19800 20204 19852 20256
rect 21456 20204 21508 20256
rect 1918 20102 1970 20154
rect 1982 20102 2034 20154
rect 2046 20102 2098 20154
rect 2110 20102 2162 20154
rect 2174 20102 2226 20154
rect 2238 20102 2290 20154
rect 7918 20102 7970 20154
rect 7982 20102 8034 20154
rect 8046 20102 8098 20154
rect 8110 20102 8162 20154
rect 8174 20102 8226 20154
rect 8238 20102 8290 20154
rect 13918 20102 13970 20154
rect 13982 20102 14034 20154
rect 14046 20102 14098 20154
rect 14110 20102 14162 20154
rect 14174 20102 14226 20154
rect 14238 20102 14290 20154
rect 19918 20102 19970 20154
rect 19982 20102 20034 20154
rect 20046 20102 20098 20154
rect 20110 20102 20162 20154
rect 20174 20102 20226 20154
rect 20238 20102 20290 20154
rect 5632 20000 5684 20052
rect 6552 20000 6604 20052
rect 9128 19864 9180 19916
rect 9496 19932 9548 19984
rect 9588 19975 9640 19984
rect 9588 19941 9597 19975
rect 9597 19941 9631 19975
rect 9631 19941 9640 19975
rect 9588 19932 9640 19941
rect 8484 19839 8536 19848
rect 8484 19805 8493 19839
rect 8493 19805 8527 19839
rect 8527 19805 8536 19839
rect 8484 19796 8536 19805
rect 8576 19796 8628 19848
rect 8668 19796 8720 19848
rect 9312 19796 9364 19848
rect 9496 19839 9548 19848
rect 9496 19805 9505 19839
rect 9505 19805 9539 19839
rect 9539 19805 9548 19839
rect 9496 19796 9548 19805
rect 9864 19796 9916 19848
rect 11612 19796 11664 19848
rect 12624 20000 12676 20052
rect 12992 20000 13044 20052
rect 14372 20000 14424 20052
rect 17776 20000 17828 20052
rect 15292 19932 15344 19984
rect 12532 19796 12584 19848
rect 13268 19796 13320 19848
rect 13820 19796 13872 19848
rect 6276 19728 6328 19780
rect 6368 19728 6420 19780
rect 7840 19728 7892 19780
rect 8300 19728 8352 19780
rect 5264 19703 5316 19712
rect 5264 19669 5273 19703
rect 5273 19669 5307 19703
rect 5307 19669 5316 19703
rect 5264 19660 5316 19669
rect 8576 19703 8628 19712
rect 8576 19669 8585 19703
rect 8585 19669 8619 19703
rect 8619 19669 8628 19703
rect 8576 19660 8628 19669
rect 10876 19728 10928 19780
rect 12072 19728 12124 19780
rect 9680 19660 9732 19712
rect 14464 19796 14516 19848
rect 15200 19839 15252 19848
rect 15200 19805 15209 19839
rect 15209 19805 15243 19839
rect 15243 19805 15252 19839
rect 15200 19796 15252 19805
rect 15476 19796 15528 19848
rect 17040 19771 17092 19780
rect 17040 19737 17049 19771
rect 17049 19737 17083 19771
rect 17083 19737 17092 19771
rect 17040 19728 17092 19737
rect 18052 19728 18104 19780
rect 18512 19839 18564 19848
rect 18512 19805 18521 19839
rect 18521 19805 18555 19839
rect 18555 19805 18564 19839
rect 18512 19796 18564 19805
rect 19340 19796 19392 19848
rect 19524 19839 19576 19848
rect 19524 19805 19558 19839
rect 19558 19805 19576 19839
rect 19524 19796 19576 19805
rect 14556 19660 14608 19712
rect 18144 19660 18196 19712
rect 18696 19703 18748 19712
rect 18696 19669 18705 19703
rect 18705 19669 18739 19703
rect 18739 19669 18748 19703
rect 18696 19660 18748 19669
rect 18972 19703 19024 19712
rect 18972 19669 18981 19703
rect 18981 19669 19015 19703
rect 19015 19669 19024 19703
rect 18972 19660 19024 19669
rect 19340 19660 19392 19712
rect 21364 19660 21416 19712
rect 2658 19558 2710 19610
rect 2722 19558 2774 19610
rect 2786 19558 2838 19610
rect 2850 19558 2902 19610
rect 2914 19558 2966 19610
rect 2978 19558 3030 19610
rect 8658 19558 8710 19610
rect 8722 19558 8774 19610
rect 8786 19558 8838 19610
rect 8850 19558 8902 19610
rect 8914 19558 8966 19610
rect 8978 19558 9030 19610
rect 14658 19558 14710 19610
rect 14722 19558 14774 19610
rect 14786 19558 14838 19610
rect 14850 19558 14902 19610
rect 14914 19558 14966 19610
rect 14978 19558 15030 19610
rect 20658 19558 20710 19610
rect 20722 19558 20774 19610
rect 20786 19558 20838 19610
rect 20850 19558 20902 19610
rect 20914 19558 20966 19610
rect 20978 19558 21030 19610
rect 5264 19456 5316 19508
rect 4620 19320 4672 19372
rect 4804 19363 4856 19372
rect 4804 19329 4813 19363
rect 4813 19329 4847 19363
rect 4847 19329 4856 19363
rect 4804 19320 4856 19329
rect 5080 19363 5132 19372
rect 5080 19329 5114 19363
rect 5114 19329 5132 19363
rect 5080 19320 5132 19329
rect 7012 19388 7064 19440
rect 7564 19456 7616 19508
rect 8392 19456 8444 19508
rect 9496 19456 9548 19508
rect 13728 19456 13780 19508
rect 14372 19456 14424 19508
rect 15200 19456 15252 19508
rect 8392 19363 8444 19372
rect 8392 19329 8426 19363
rect 8426 19329 8444 19363
rect 8392 19320 8444 19329
rect 9220 19320 9272 19372
rect 10140 19320 10192 19372
rect 10692 19320 10744 19372
rect 10784 19252 10836 19304
rect 11060 19252 11112 19304
rect 11704 19363 11756 19372
rect 11704 19329 11713 19363
rect 11713 19329 11747 19363
rect 11747 19329 11756 19363
rect 11704 19320 11756 19329
rect 11888 19252 11940 19304
rect 21364 19456 21416 19508
rect 13176 19320 13228 19372
rect 14372 19320 14424 19372
rect 16764 19388 16816 19440
rect 17408 19388 17460 19440
rect 15108 19320 15160 19372
rect 14556 19295 14608 19304
rect 14556 19261 14565 19295
rect 14565 19261 14599 19295
rect 14599 19261 14608 19295
rect 14556 19252 14608 19261
rect 17224 19320 17276 19372
rect 18144 19320 18196 19372
rect 19524 19388 19576 19440
rect 18420 19320 18472 19372
rect 19340 19320 19392 19372
rect 23296 19363 23348 19372
rect 23296 19329 23305 19363
rect 23305 19329 23339 19363
rect 23339 19329 23348 19363
rect 23296 19320 23348 19329
rect 18236 19295 18288 19304
rect 18236 19261 18245 19295
rect 18245 19261 18279 19295
rect 18279 19261 18288 19295
rect 18236 19252 18288 19261
rect 4528 19159 4580 19168
rect 4528 19125 4537 19159
rect 4537 19125 4571 19159
rect 4571 19125 4580 19159
rect 4528 19116 4580 19125
rect 5908 19116 5960 19168
rect 9772 19116 9824 19168
rect 10876 19116 10928 19168
rect 16672 19184 16724 19236
rect 14924 19116 14976 19168
rect 20444 19295 20496 19304
rect 20444 19261 20453 19295
rect 20453 19261 20487 19295
rect 20487 19261 20496 19295
rect 20444 19252 20496 19261
rect 19616 19184 19668 19236
rect 19708 19159 19760 19168
rect 19708 19125 19717 19159
rect 19717 19125 19751 19159
rect 19751 19125 19760 19159
rect 19708 19116 19760 19125
rect 1918 19014 1970 19066
rect 1982 19014 2034 19066
rect 2046 19014 2098 19066
rect 2110 19014 2162 19066
rect 2174 19014 2226 19066
rect 2238 19014 2290 19066
rect 7918 19014 7970 19066
rect 7982 19014 8034 19066
rect 8046 19014 8098 19066
rect 8110 19014 8162 19066
rect 8174 19014 8226 19066
rect 8238 19014 8290 19066
rect 13918 19014 13970 19066
rect 13982 19014 14034 19066
rect 14046 19014 14098 19066
rect 14110 19014 14162 19066
rect 14174 19014 14226 19066
rect 14238 19014 14290 19066
rect 19918 19014 19970 19066
rect 19982 19014 20034 19066
rect 20046 19014 20098 19066
rect 20110 19014 20162 19066
rect 20174 19014 20226 19066
rect 20238 19014 20290 19066
rect 5080 18912 5132 18964
rect 6736 18955 6788 18964
rect 6736 18921 6745 18955
rect 6745 18921 6779 18955
rect 6779 18921 6788 18955
rect 6736 18912 6788 18921
rect 9864 18912 9916 18964
rect 10048 18912 10100 18964
rect 14556 18912 14608 18964
rect 18236 18912 18288 18964
rect 20444 18912 20496 18964
rect 9588 18844 9640 18896
rect 6828 18819 6880 18828
rect 6828 18785 6837 18819
rect 6837 18785 6871 18819
rect 6871 18785 6880 18819
rect 6828 18776 6880 18785
rect 3884 18751 3936 18760
rect 3884 18717 3893 18751
rect 3893 18717 3927 18751
rect 3927 18717 3936 18751
rect 3884 18708 3936 18717
rect 4528 18708 4580 18760
rect 5356 18751 5408 18760
rect 5356 18717 5365 18751
rect 5365 18717 5399 18751
rect 5399 18717 5408 18751
rect 5356 18708 5408 18717
rect 5908 18708 5960 18760
rect 6920 18708 6972 18760
rect 4620 18640 4672 18692
rect 5540 18640 5592 18692
rect 11520 18776 11572 18828
rect 15476 18844 15528 18896
rect 8484 18708 8536 18760
rect 10508 18751 10560 18760
rect 10508 18717 10517 18751
rect 10517 18717 10551 18751
rect 10551 18717 10560 18751
rect 10508 18708 10560 18717
rect 10968 18751 11020 18760
rect 10968 18717 10977 18751
rect 10977 18717 11011 18751
rect 11011 18717 11020 18751
rect 10968 18708 11020 18717
rect 11152 18751 11204 18760
rect 11152 18717 11161 18751
rect 11161 18717 11195 18751
rect 11195 18717 11204 18751
rect 11152 18708 11204 18717
rect 9496 18640 9548 18692
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 14648 18776 14700 18828
rect 15200 18776 15252 18828
rect 14464 18708 14516 18760
rect 14556 18708 14608 18760
rect 18696 18776 18748 18828
rect 18972 18776 19024 18828
rect 18880 18751 18932 18760
rect 18880 18717 18889 18751
rect 18889 18717 18923 18751
rect 18923 18717 18932 18751
rect 18880 18708 18932 18717
rect 10048 18572 10100 18624
rect 11428 18572 11480 18624
rect 11796 18572 11848 18624
rect 11980 18572 12032 18624
rect 13820 18640 13872 18692
rect 14004 18640 14056 18692
rect 21272 18751 21324 18760
rect 21272 18717 21281 18751
rect 21281 18717 21315 18751
rect 21315 18717 21324 18751
rect 21272 18708 21324 18717
rect 21456 18708 21508 18760
rect 19800 18640 19852 18692
rect 23296 18683 23348 18692
rect 23296 18649 23305 18683
rect 23305 18649 23339 18683
rect 23339 18649 23348 18683
rect 23296 18640 23348 18649
rect 13176 18615 13228 18624
rect 13176 18581 13185 18615
rect 13185 18581 13219 18615
rect 13219 18581 13228 18615
rect 13176 18572 13228 18581
rect 13544 18572 13596 18624
rect 14280 18572 14332 18624
rect 17960 18615 18012 18624
rect 17960 18581 17969 18615
rect 17969 18581 18003 18615
rect 18003 18581 18012 18615
rect 17960 18572 18012 18581
rect 2658 18470 2710 18522
rect 2722 18470 2774 18522
rect 2786 18470 2838 18522
rect 2850 18470 2902 18522
rect 2914 18470 2966 18522
rect 2978 18470 3030 18522
rect 8658 18470 8710 18522
rect 8722 18470 8774 18522
rect 8786 18470 8838 18522
rect 8850 18470 8902 18522
rect 8914 18470 8966 18522
rect 8978 18470 9030 18522
rect 14658 18470 14710 18522
rect 14722 18470 14774 18522
rect 14786 18470 14838 18522
rect 14850 18470 14902 18522
rect 14914 18470 14966 18522
rect 14978 18470 15030 18522
rect 20658 18470 20710 18522
rect 20722 18470 20774 18522
rect 20786 18470 20838 18522
rect 20850 18470 20902 18522
rect 20914 18470 20966 18522
rect 20978 18470 21030 18522
rect 3884 18368 3936 18420
rect 5356 18368 5408 18420
rect 5448 18368 5500 18420
rect 4160 18275 4212 18284
rect 4160 18241 4169 18275
rect 4169 18241 4203 18275
rect 4203 18241 4212 18275
rect 4160 18232 4212 18241
rect 6276 18300 6328 18352
rect 9312 18368 9364 18420
rect 10048 18368 10100 18420
rect 14004 18368 14056 18420
rect 14372 18368 14424 18420
rect 15108 18368 15160 18420
rect 18052 18411 18104 18420
rect 18052 18377 18061 18411
rect 18061 18377 18095 18411
rect 18095 18377 18104 18411
rect 18052 18368 18104 18377
rect 18144 18411 18196 18420
rect 18144 18377 18153 18411
rect 18153 18377 18187 18411
rect 18187 18377 18196 18411
rect 18144 18368 18196 18377
rect 21272 18368 21324 18420
rect 16856 18300 16908 18352
rect 19708 18300 19760 18352
rect 5540 18232 5592 18284
rect 6092 18232 6144 18284
rect 6184 18275 6236 18284
rect 6184 18241 6193 18275
rect 6193 18241 6227 18275
rect 6227 18241 6236 18275
rect 6184 18232 6236 18241
rect 6736 18232 6788 18284
rect 7472 18232 7524 18284
rect 10600 18232 10652 18284
rect 14464 18232 14516 18284
rect 16764 18232 16816 18284
rect 16948 18275 17000 18284
rect 16948 18241 16982 18275
rect 16982 18241 17000 18275
rect 16948 18232 17000 18241
rect 4896 18164 4948 18216
rect 9864 18164 9916 18216
rect 11888 18164 11940 18216
rect 13268 18164 13320 18216
rect 19524 18207 19576 18216
rect 19524 18173 19533 18207
rect 19533 18173 19567 18207
rect 19567 18173 19576 18207
rect 19524 18164 19576 18173
rect 19616 18207 19668 18216
rect 19616 18173 19625 18207
rect 19625 18173 19659 18207
rect 19659 18173 19668 18207
rect 19616 18164 19668 18173
rect 7840 18096 7892 18148
rect 11244 18096 11296 18148
rect 14648 18096 14700 18148
rect 15200 18096 15252 18148
rect 4896 18028 4948 18080
rect 6276 18028 6328 18080
rect 8392 18028 8444 18080
rect 14740 18028 14792 18080
rect 1918 17926 1970 17978
rect 1982 17926 2034 17978
rect 2046 17926 2098 17978
rect 2110 17926 2162 17978
rect 2174 17926 2226 17978
rect 2238 17926 2290 17978
rect 7918 17926 7970 17978
rect 7982 17926 8034 17978
rect 8046 17926 8098 17978
rect 8110 17926 8162 17978
rect 8174 17926 8226 17978
rect 8238 17926 8290 17978
rect 13918 17926 13970 17978
rect 13982 17926 14034 17978
rect 14046 17926 14098 17978
rect 14110 17926 14162 17978
rect 14174 17926 14226 17978
rect 14238 17926 14290 17978
rect 19918 17926 19970 17978
rect 19982 17926 20034 17978
rect 20046 17926 20098 17978
rect 20110 17926 20162 17978
rect 20174 17926 20226 17978
rect 20238 17926 20290 17978
rect 7472 17824 7524 17876
rect 10600 17824 10652 17876
rect 11152 17824 11204 17876
rect 13360 17824 13412 17876
rect 14648 17824 14700 17876
rect 4712 17756 4764 17808
rect 4252 17688 4304 17740
rect 7012 17731 7064 17740
rect 7012 17697 7021 17731
rect 7021 17697 7055 17731
rect 7055 17697 7064 17731
rect 7012 17688 7064 17697
rect 5356 17620 5408 17672
rect 3516 17484 3568 17536
rect 4160 17484 4212 17536
rect 6552 17595 6604 17604
rect 6552 17561 6561 17595
rect 6561 17561 6595 17595
rect 6595 17561 6604 17595
rect 6552 17552 6604 17561
rect 8484 17552 8536 17604
rect 11612 17799 11664 17808
rect 11612 17765 11621 17799
rect 11621 17765 11655 17799
rect 11655 17765 11664 17799
rect 11612 17756 11664 17765
rect 16948 17824 17000 17876
rect 18512 17824 18564 17876
rect 17960 17756 18012 17808
rect 18880 17756 18932 17808
rect 9680 17688 9732 17740
rect 9128 17620 9180 17672
rect 11704 17688 11756 17740
rect 11888 17620 11940 17672
rect 10692 17552 10744 17604
rect 12072 17552 12124 17604
rect 13728 17663 13780 17672
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 13728 17620 13780 17629
rect 14372 17620 14424 17672
rect 18052 17620 18104 17672
rect 19064 17620 19116 17672
rect 19340 17663 19392 17672
rect 19340 17629 19349 17663
rect 19349 17629 19383 17663
rect 19383 17629 19392 17663
rect 19340 17620 19392 17629
rect 15108 17552 15160 17604
rect 6828 17527 6880 17536
rect 6828 17493 6837 17527
rect 6837 17493 6871 17527
rect 6871 17493 6880 17527
rect 6828 17484 6880 17493
rect 6920 17484 6972 17536
rect 13636 17527 13688 17536
rect 13636 17493 13645 17527
rect 13645 17493 13679 17527
rect 13679 17493 13688 17527
rect 13636 17484 13688 17493
rect 14372 17484 14424 17536
rect 14740 17484 14792 17536
rect 16488 17484 16540 17536
rect 18144 17527 18196 17536
rect 18144 17493 18153 17527
rect 18153 17493 18187 17527
rect 18187 17493 18196 17527
rect 18144 17484 18196 17493
rect 18972 17527 19024 17536
rect 18972 17493 18981 17527
rect 18981 17493 19015 17527
rect 19015 17493 19024 17527
rect 18972 17484 19024 17493
rect 19432 17527 19484 17536
rect 19432 17493 19441 17527
rect 19441 17493 19475 17527
rect 19475 17493 19484 17527
rect 19432 17484 19484 17493
rect 2658 17382 2710 17434
rect 2722 17382 2774 17434
rect 2786 17382 2838 17434
rect 2850 17382 2902 17434
rect 2914 17382 2966 17434
rect 2978 17382 3030 17434
rect 8658 17382 8710 17434
rect 8722 17382 8774 17434
rect 8786 17382 8838 17434
rect 8850 17382 8902 17434
rect 8914 17382 8966 17434
rect 8978 17382 9030 17434
rect 14658 17382 14710 17434
rect 14722 17382 14774 17434
rect 14786 17382 14838 17434
rect 14850 17382 14902 17434
rect 14914 17382 14966 17434
rect 14978 17382 15030 17434
rect 20658 17382 20710 17434
rect 20722 17382 20774 17434
rect 20786 17382 20838 17434
rect 20850 17382 20902 17434
rect 20914 17382 20966 17434
rect 20978 17382 21030 17434
rect 4712 17323 4764 17332
rect 4712 17289 4721 17323
rect 4721 17289 4755 17323
rect 4755 17289 4764 17323
rect 4712 17280 4764 17289
rect 6552 17280 6604 17332
rect 6736 17323 6788 17332
rect 6736 17289 6745 17323
rect 6745 17289 6779 17323
rect 6779 17289 6788 17323
rect 6736 17280 6788 17289
rect 6920 17280 6972 17332
rect 3332 17144 3384 17196
rect 3424 17187 3476 17196
rect 3424 17153 3433 17187
rect 3433 17153 3467 17187
rect 3467 17153 3476 17187
rect 3424 17144 3476 17153
rect 4528 17212 4580 17264
rect 3976 17187 4028 17196
rect 3976 17153 3985 17187
rect 3985 17153 4019 17187
rect 4019 17153 4028 17187
rect 3976 17144 4028 17153
rect 4252 17144 4304 17196
rect 4436 17144 4488 17196
rect 4804 17187 4856 17196
rect 4804 17153 4813 17187
rect 4813 17153 4847 17187
rect 4847 17153 4856 17187
rect 4804 17144 4856 17153
rect 940 17076 992 17128
rect 6368 17212 6420 17264
rect 5080 17187 5132 17196
rect 5080 17153 5114 17187
rect 5114 17153 5132 17187
rect 5080 17144 5132 17153
rect 4620 17008 4672 17060
rect 3056 16940 3108 16992
rect 4252 16940 4304 16992
rect 5172 16940 5224 16992
rect 7104 17076 7156 17128
rect 9404 17280 9456 17332
rect 13268 17323 13320 17332
rect 13268 17289 13277 17323
rect 13277 17289 13311 17323
rect 13311 17289 13320 17323
rect 13268 17280 13320 17289
rect 13636 17280 13688 17332
rect 15660 17280 15712 17332
rect 16856 17280 16908 17332
rect 17040 17280 17092 17332
rect 17868 17280 17920 17332
rect 18144 17280 18196 17332
rect 18972 17280 19024 17332
rect 13176 17212 13228 17264
rect 11428 17144 11480 17196
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 14372 17212 14424 17264
rect 15292 17187 15344 17196
rect 15292 17153 15326 17187
rect 15326 17153 15344 17187
rect 15292 17144 15344 17153
rect 16856 17144 16908 17196
rect 19616 17187 19668 17196
rect 19616 17153 19634 17187
rect 19634 17153 19668 17187
rect 19616 17144 19668 17153
rect 21180 17144 21232 17196
rect 7012 17008 7064 17060
rect 11520 17008 11572 17060
rect 5908 16940 5960 16992
rect 6460 16940 6512 16992
rect 10508 16940 10560 16992
rect 18512 16983 18564 16992
rect 18512 16949 18521 16983
rect 18521 16949 18555 16983
rect 18555 16949 18564 16983
rect 18512 16940 18564 16949
rect 19524 16940 19576 16992
rect 23296 17119 23348 17128
rect 23296 17085 23305 17119
rect 23305 17085 23339 17119
rect 23339 17085 23348 17119
rect 23296 17076 23348 17085
rect 21088 16940 21140 16992
rect 1918 16838 1970 16890
rect 1982 16838 2034 16890
rect 2046 16838 2098 16890
rect 2110 16838 2162 16890
rect 2174 16838 2226 16890
rect 2238 16838 2290 16890
rect 7918 16838 7970 16890
rect 7982 16838 8034 16890
rect 8046 16838 8098 16890
rect 8110 16838 8162 16890
rect 8174 16838 8226 16890
rect 8238 16838 8290 16890
rect 13918 16838 13970 16890
rect 13982 16838 14034 16890
rect 14046 16838 14098 16890
rect 14110 16838 14162 16890
rect 14174 16838 14226 16890
rect 14238 16838 14290 16890
rect 19918 16838 19970 16890
rect 19982 16838 20034 16890
rect 20046 16838 20098 16890
rect 20110 16838 20162 16890
rect 20174 16838 20226 16890
rect 20238 16838 20290 16890
rect 6092 16736 6144 16788
rect 6184 16736 6236 16788
rect 6828 16736 6880 16788
rect 11612 16779 11664 16788
rect 11612 16745 11621 16779
rect 11621 16745 11655 16779
rect 11655 16745 11664 16779
rect 11612 16736 11664 16745
rect 18420 16736 18472 16788
rect 19892 16736 19944 16788
rect 21180 16779 21232 16788
rect 21180 16745 21189 16779
rect 21189 16745 21223 16779
rect 21223 16745 21232 16779
rect 21180 16736 21232 16745
rect 3240 16600 3292 16652
rect 2136 16575 2188 16584
rect 2136 16541 2145 16575
rect 2145 16541 2179 16575
rect 2179 16541 2188 16575
rect 2136 16532 2188 16541
rect 5172 16600 5224 16652
rect 9036 16711 9088 16720
rect 9036 16677 9045 16711
rect 9045 16677 9079 16711
rect 9079 16677 9088 16711
rect 9036 16668 9088 16677
rect 5816 16532 5868 16584
rect 6276 16532 6328 16584
rect 14372 16600 14424 16652
rect 18052 16600 18104 16652
rect 19800 16668 19852 16720
rect 21732 16668 21784 16720
rect 4160 16464 4212 16516
rect 15844 16575 15896 16584
rect 1216 16396 1268 16448
rect 2412 16396 2464 16448
rect 3424 16396 3476 16448
rect 4068 16439 4120 16448
rect 4068 16405 4077 16439
rect 4077 16405 4111 16439
rect 4111 16405 4120 16439
rect 4068 16396 4120 16405
rect 5448 16396 5500 16448
rect 8668 16464 8720 16516
rect 9404 16507 9456 16516
rect 9404 16473 9413 16507
rect 9413 16473 9447 16507
rect 9447 16473 9456 16507
rect 9404 16464 9456 16473
rect 7748 16396 7800 16448
rect 8300 16439 8352 16448
rect 8300 16405 8309 16439
rect 8309 16405 8343 16439
rect 8343 16405 8352 16439
rect 8300 16396 8352 16405
rect 9864 16439 9916 16448
rect 9864 16405 9873 16439
rect 9873 16405 9907 16439
rect 9907 16405 9916 16439
rect 9864 16396 9916 16405
rect 13544 16464 13596 16516
rect 13176 16396 13228 16448
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 18420 16575 18472 16584
rect 18420 16541 18429 16575
rect 18429 16541 18463 16575
rect 18463 16541 18472 16575
rect 18420 16532 18472 16541
rect 21088 16643 21140 16652
rect 21088 16609 21097 16643
rect 21097 16609 21131 16643
rect 21131 16609 21140 16643
rect 21088 16600 21140 16609
rect 22192 16600 22244 16652
rect 15936 16507 15988 16516
rect 15936 16473 15945 16507
rect 15945 16473 15979 16507
rect 15979 16473 15988 16507
rect 15936 16464 15988 16473
rect 18604 16464 18656 16516
rect 23020 16575 23072 16584
rect 23020 16541 23029 16575
rect 23029 16541 23063 16575
rect 23063 16541 23072 16575
rect 23020 16532 23072 16541
rect 23204 16464 23256 16516
rect 13820 16396 13872 16448
rect 16212 16396 16264 16448
rect 18236 16396 18288 16448
rect 19248 16396 19300 16448
rect 19340 16439 19392 16448
rect 19340 16405 19349 16439
rect 19349 16405 19383 16439
rect 19383 16405 19392 16439
rect 19340 16396 19392 16405
rect 19708 16439 19760 16448
rect 19708 16405 19717 16439
rect 19717 16405 19751 16439
rect 19751 16405 19760 16439
rect 19708 16396 19760 16405
rect 21916 16439 21968 16448
rect 21916 16405 21925 16439
rect 21925 16405 21959 16439
rect 21959 16405 21968 16439
rect 21916 16396 21968 16405
rect 22744 16439 22796 16448
rect 22744 16405 22753 16439
rect 22753 16405 22787 16439
rect 22787 16405 22796 16439
rect 22744 16396 22796 16405
rect 23112 16396 23164 16448
rect 2658 16294 2710 16346
rect 2722 16294 2774 16346
rect 2786 16294 2838 16346
rect 2850 16294 2902 16346
rect 2914 16294 2966 16346
rect 2978 16294 3030 16346
rect 8658 16294 8710 16346
rect 8722 16294 8774 16346
rect 8786 16294 8838 16346
rect 8850 16294 8902 16346
rect 8914 16294 8966 16346
rect 8978 16294 9030 16346
rect 14658 16294 14710 16346
rect 14722 16294 14774 16346
rect 14786 16294 14838 16346
rect 14850 16294 14902 16346
rect 14914 16294 14966 16346
rect 14978 16294 15030 16346
rect 20658 16294 20710 16346
rect 20722 16294 20774 16346
rect 20786 16294 20838 16346
rect 20850 16294 20902 16346
rect 20914 16294 20966 16346
rect 20978 16294 21030 16346
rect 3332 16235 3384 16244
rect 3332 16201 3341 16235
rect 3341 16201 3375 16235
rect 3375 16201 3384 16235
rect 3332 16192 3384 16201
rect 3700 16192 3752 16244
rect 9772 16192 9824 16244
rect 11520 16235 11572 16244
rect 11520 16201 11529 16235
rect 11529 16201 11563 16235
rect 11563 16201 11572 16235
rect 11520 16192 11572 16201
rect 12072 16235 12124 16244
rect 12072 16201 12081 16235
rect 12081 16201 12115 16235
rect 12115 16201 12124 16235
rect 12072 16192 12124 16201
rect 1492 16124 1544 16176
rect 1860 16099 1912 16108
rect 1860 16065 1869 16099
rect 1869 16065 1903 16099
rect 1903 16065 1912 16099
rect 1860 16056 1912 16065
rect 3424 16124 3476 16176
rect 940 15988 992 16040
rect 1676 15988 1728 16040
rect 2504 15988 2556 16040
rect 3700 16056 3752 16108
rect 4068 16124 4120 16176
rect 4896 16124 4948 16176
rect 6644 16099 6696 16108
rect 6644 16065 6653 16099
rect 6653 16065 6687 16099
rect 6687 16065 6696 16099
rect 6644 16056 6696 16065
rect 7012 16056 7064 16108
rect 7840 16099 7892 16108
rect 11888 16124 11940 16176
rect 13268 16192 13320 16244
rect 14372 16235 14424 16244
rect 14372 16201 14381 16235
rect 14381 16201 14415 16235
rect 14415 16201 14424 16235
rect 14372 16192 14424 16201
rect 15844 16192 15896 16244
rect 13912 16124 13964 16176
rect 17040 16192 17092 16244
rect 19524 16192 19576 16244
rect 19800 16192 19852 16244
rect 7840 16065 7858 16099
rect 7858 16065 7892 16099
rect 7840 16056 7892 16065
rect 3608 15988 3660 16040
rect 4712 16031 4764 16040
rect 4712 15997 4721 16031
rect 4721 15997 4755 16031
rect 4755 15997 4764 16031
rect 4712 15988 4764 15997
rect 2504 15895 2556 15904
rect 2504 15861 2513 15895
rect 2513 15861 2547 15895
rect 2547 15861 2556 15895
rect 2504 15852 2556 15861
rect 3700 15852 3752 15904
rect 4528 15852 4580 15904
rect 7012 15920 7064 15972
rect 6368 15852 6420 15904
rect 6828 15852 6880 15904
rect 13820 16056 13872 16108
rect 11336 16031 11388 16040
rect 11336 15997 11345 16031
rect 11345 15997 11379 16031
rect 11379 15997 11388 16031
rect 11336 15988 11388 15997
rect 13728 15988 13780 16040
rect 14372 16056 14424 16108
rect 14556 16056 14608 16108
rect 15292 16056 15344 16108
rect 17868 16124 17920 16176
rect 9496 15963 9548 15972
rect 9496 15929 9505 15963
rect 9505 15929 9539 15963
rect 9539 15929 9548 15963
rect 9496 15920 9548 15929
rect 11796 15920 11848 15972
rect 9680 15852 9732 15904
rect 13452 15852 13504 15904
rect 16672 16099 16724 16108
rect 16672 16065 16681 16099
rect 16681 16065 16715 16099
rect 16715 16065 16724 16099
rect 16672 16056 16724 16065
rect 23112 16124 23164 16176
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 20352 15988 20404 16040
rect 22100 16031 22152 16040
rect 22100 15997 22109 16031
rect 22109 15997 22143 16031
rect 22143 15997 22152 16031
rect 22100 15988 22152 15997
rect 22928 15988 22980 16040
rect 19064 15920 19116 15972
rect 21640 15920 21692 15972
rect 23204 15920 23256 15972
rect 15108 15852 15160 15904
rect 16120 15895 16172 15904
rect 16120 15861 16129 15895
rect 16129 15861 16163 15895
rect 16163 15861 16172 15895
rect 16120 15852 16172 15861
rect 16580 15852 16632 15904
rect 17960 15852 18012 15904
rect 21456 15895 21508 15904
rect 21456 15861 21465 15895
rect 21465 15861 21499 15895
rect 21499 15861 21508 15895
rect 21456 15852 21508 15861
rect 22560 15852 22612 15904
rect 22836 15895 22888 15904
rect 22836 15861 22845 15895
rect 22845 15861 22879 15895
rect 22879 15861 22888 15895
rect 22836 15852 22888 15861
rect 1918 15750 1970 15802
rect 1982 15750 2034 15802
rect 2046 15750 2098 15802
rect 2110 15750 2162 15802
rect 2174 15750 2226 15802
rect 2238 15750 2290 15802
rect 7918 15750 7970 15802
rect 7982 15750 8034 15802
rect 8046 15750 8098 15802
rect 8110 15750 8162 15802
rect 8174 15750 8226 15802
rect 8238 15750 8290 15802
rect 13918 15750 13970 15802
rect 13982 15750 14034 15802
rect 14046 15750 14098 15802
rect 14110 15750 14162 15802
rect 14174 15750 14226 15802
rect 14238 15750 14290 15802
rect 19918 15750 19970 15802
rect 19982 15750 20034 15802
rect 20046 15750 20098 15802
rect 20110 15750 20162 15802
rect 20174 15750 20226 15802
rect 20238 15750 20290 15802
rect 3884 15648 3936 15700
rect 4712 15648 4764 15700
rect 4804 15648 4856 15700
rect 7472 15648 7524 15700
rect 8576 15648 8628 15700
rect 4068 15580 4120 15632
rect 5448 15580 5500 15632
rect 2228 15444 2280 15496
rect 3516 15512 3568 15564
rect 4252 15512 4304 15564
rect 11980 15691 12032 15700
rect 11980 15657 11989 15691
rect 11989 15657 12023 15691
rect 12023 15657 12032 15691
rect 11980 15648 12032 15657
rect 13728 15648 13780 15700
rect 15384 15648 15436 15700
rect 15476 15648 15528 15700
rect 16120 15648 16172 15700
rect 17132 15648 17184 15700
rect 17040 15580 17092 15632
rect 10508 15512 10560 15564
rect 1860 15376 1912 15428
rect 1584 15308 1636 15360
rect 1768 15308 1820 15360
rect 2136 15351 2188 15360
rect 2136 15317 2145 15351
rect 2145 15317 2179 15351
rect 2179 15317 2188 15351
rect 2136 15308 2188 15317
rect 2412 15308 2464 15360
rect 3608 15444 3660 15496
rect 3700 15444 3752 15496
rect 3976 15444 4028 15496
rect 4528 15444 4580 15496
rect 3332 15308 3384 15360
rect 9864 15444 9916 15496
rect 10876 15487 10928 15496
rect 10876 15453 10910 15487
rect 10910 15453 10928 15487
rect 10876 15444 10928 15453
rect 12072 15487 12124 15496
rect 12072 15453 12081 15487
rect 12081 15453 12115 15487
rect 12115 15453 12124 15487
rect 12072 15444 12124 15453
rect 14372 15512 14424 15564
rect 16488 15512 16540 15564
rect 16948 15512 17000 15564
rect 19340 15648 19392 15700
rect 18880 15580 18932 15632
rect 21088 15580 21140 15632
rect 17592 15487 17644 15496
rect 17592 15453 17601 15487
rect 17601 15453 17635 15487
rect 17635 15453 17644 15487
rect 17592 15444 17644 15453
rect 22560 15444 22612 15496
rect 22652 15444 22704 15496
rect 4712 15419 4764 15428
rect 4712 15385 4746 15419
rect 4746 15385 4764 15419
rect 4712 15376 4764 15385
rect 8392 15376 8444 15428
rect 9956 15376 10008 15428
rect 12348 15419 12400 15428
rect 12348 15385 12382 15419
rect 12382 15385 12400 15419
rect 12348 15376 12400 15385
rect 15200 15376 15252 15428
rect 15476 15419 15528 15428
rect 15476 15385 15516 15419
rect 15516 15385 15528 15419
rect 15476 15376 15528 15385
rect 9220 15308 9272 15360
rect 13820 15351 13872 15360
rect 13820 15317 13829 15351
rect 13829 15317 13863 15351
rect 13863 15317 13872 15351
rect 13820 15308 13872 15317
rect 14556 15308 14608 15360
rect 18144 15376 18196 15428
rect 19524 15376 19576 15428
rect 23020 15376 23072 15428
rect 19616 15308 19668 15360
rect 21364 15308 21416 15360
rect 22560 15351 22612 15360
rect 22560 15317 22569 15351
rect 22569 15317 22603 15351
rect 22603 15317 22612 15351
rect 22560 15308 22612 15317
rect 23112 15308 23164 15360
rect 2658 15206 2710 15258
rect 2722 15206 2774 15258
rect 2786 15206 2838 15258
rect 2850 15206 2902 15258
rect 2914 15206 2966 15258
rect 2978 15206 3030 15258
rect 8658 15206 8710 15258
rect 8722 15206 8774 15258
rect 8786 15206 8838 15258
rect 8850 15206 8902 15258
rect 8914 15206 8966 15258
rect 8978 15206 9030 15258
rect 14658 15206 14710 15258
rect 14722 15206 14774 15258
rect 14786 15206 14838 15258
rect 14850 15206 14902 15258
rect 14914 15206 14966 15258
rect 14978 15206 15030 15258
rect 20658 15206 20710 15258
rect 20722 15206 20774 15258
rect 20786 15206 20838 15258
rect 20850 15206 20902 15258
rect 20914 15206 20966 15258
rect 20978 15206 21030 15258
rect 1584 15104 1636 15156
rect 3240 15104 3292 15156
rect 3056 15036 3108 15088
rect 3148 14968 3200 15020
rect 4436 15104 4488 15156
rect 3700 15036 3752 15088
rect 5080 15104 5132 15156
rect 6092 15104 6144 15156
rect 7104 15104 7156 15156
rect 8484 15104 8536 15156
rect 12072 15104 12124 15156
rect 4620 15036 4672 15088
rect 1860 14943 1912 14952
rect 1860 14909 1869 14943
rect 1869 14909 1903 14943
rect 1903 14909 1912 14943
rect 1860 14900 1912 14909
rect 4160 14968 4212 15020
rect 9588 15011 9640 15020
rect 9588 14977 9597 15011
rect 9597 14977 9631 15011
rect 9631 14977 9640 15011
rect 9588 14968 9640 14977
rect 11060 15036 11112 15088
rect 9772 14968 9824 15020
rect 10784 14968 10836 15020
rect 14372 15147 14424 15156
rect 14372 15113 14381 15147
rect 14381 15113 14415 15147
rect 14415 15113 14424 15147
rect 14372 15104 14424 15113
rect 13452 15079 13504 15088
rect 13452 15045 13492 15079
rect 13492 15045 13504 15079
rect 13452 15036 13504 15045
rect 17592 15036 17644 15088
rect 19248 15036 19300 15088
rect 19708 15036 19760 15088
rect 13820 14968 13872 15020
rect 16580 14968 16632 15020
rect 17224 14968 17276 15020
rect 17684 14968 17736 15020
rect 17960 14968 18012 15020
rect 1676 14807 1728 14816
rect 1676 14773 1685 14807
rect 1685 14773 1719 14807
rect 1719 14773 1728 14807
rect 1676 14764 1728 14773
rect 2136 14764 2188 14816
rect 2596 14764 2648 14816
rect 3608 14764 3660 14816
rect 16304 14943 16356 14952
rect 16304 14909 16313 14943
rect 16313 14909 16347 14943
rect 16347 14909 16356 14943
rect 16304 14900 16356 14909
rect 19432 14968 19484 15020
rect 21088 15104 21140 15156
rect 22100 15104 22152 15156
rect 21640 15036 21692 15088
rect 6368 14764 6420 14816
rect 9956 14764 10008 14816
rect 10968 14764 11020 14816
rect 11336 14807 11388 14816
rect 11336 14773 11345 14807
rect 11345 14773 11379 14807
rect 11379 14773 11388 14807
rect 11336 14764 11388 14773
rect 11612 14807 11664 14816
rect 11612 14773 11621 14807
rect 11621 14773 11655 14807
rect 11655 14773 11664 14807
rect 11612 14764 11664 14773
rect 14372 14764 14424 14816
rect 15752 14807 15804 14816
rect 15752 14773 15761 14807
rect 15761 14773 15795 14807
rect 15795 14773 15804 14807
rect 15752 14764 15804 14773
rect 16488 14764 16540 14816
rect 19524 14900 19576 14952
rect 20628 14900 20680 14952
rect 22376 14968 22428 15020
rect 23204 15011 23256 15020
rect 23204 14977 23213 15011
rect 23213 14977 23247 15011
rect 23247 14977 23256 15011
rect 23204 14968 23256 14977
rect 23296 15011 23348 15020
rect 23296 14977 23305 15011
rect 23305 14977 23339 15011
rect 23339 14977 23348 15011
rect 23296 14968 23348 14977
rect 19800 14764 19852 14816
rect 20536 14764 20588 14816
rect 21272 14764 21324 14816
rect 23204 14832 23256 14884
rect 22284 14764 22336 14816
rect 22468 14764 22520 14816
rect 1918 14662 1970 14714
rect 1982 14662 2034 14714
rect 2046 14662 2098 14714
rect 2110 14662 2162 14714
rect 2174 14662 2226 14714
rect 2238 14662 2290 14714
rect 7918 14662 7970 14714
rect 7982 14662 8034 14714
rect 8046 14662 8098 14714
rect 8110 14662 8162 14714
rect 8174 14662 8226 14714
rect 8238 14662 8290 14714
rect 13918 14662 13970 14714
rect 13982 14662 14034 14714
rect 14046 14662 14098 14714
rect 14110 14662 14162 14714
rect 14174 14662 14226 14714
rect 14238 14662 14290 14714
rect 19918 14662 19970 14714
rect 19982 14662 20034 14714
rect 20046 14662 20098 14714
rect 20110 14662 20162 14714
rect 20174 14662 20226 14714
rect 20238 14662 20290 14714
rect 1676 14560 1728 14612
rect 3516 14492 3568 14544
rect 3608 14535 3660 14544
rect 3608 14501 3617 14535
rect 3617 14501 3651 14535
rect 3651 14501 3660 14535
rect 3608 14492 3660 14501
rect 5080 14492 5132 14544
rect 3332 14424 3384 14476
rect 1308 14288 1360 14340
rect 2136 14288 2188 14340
rect 2596 14288 2648 14340
rect 9680 14560 9732 14612
rect 11980 14560 12032 14612
rect 16304 14560 16356 14612
rect 17040 14603 17092 14612
rect 17040 14569 17049 14603
rect 17049 14569 17083 14603
rect 17083 14569 17092 14603
rect 17040 14560 17092 14569
rect 6460 14399 6512 14408
rect 6460 14365 6478 14399
rect 6478 14365 6512 14399
rect 6460 14356 6512 14365
rect 9772 14356 9824 14408
rect 13820 14492 13872 14544
rect 15200 14424 15252 14476
rect 20536 14560 20588 14612
rect 18604 14424 18656 14476
rect 13360 14399 13412 14408
rect 13360 14365 13369 14399
rect 13369 14365 13403 14399
rect 13403 14365 13412 14399
rect 13360 14356 13412 14365
rect 15384 14356 15436 14408
rect 17132 14356 17184 14408
rect 3424 14288 3476 14340
rect 3884 14288 3936 14340
rect 4436 14288 4488 14340
rect 4712 14288 4764 14340
rect 3700 14220 3752 14272
rect 9956 14331 10008 14340
rect 9956 14297 9990 14331
rect 9990 14297 10008 14331
rect 9956 14288 10008 14297
rect 7104 14263 7156 14272
rect 7104 14229 7113 14263
rect 7113 14229 7147 14263
rect 7147 14229 7156 14263
rect 7104 14220 7156 14229
rect 7288 14220 7340 14272
rect 9496 14220 9548 14272
rect 12164 14288 12216 14340
rect 14188 14288 14240 14340
rect 11152 14220 11204 14272
rect 13544 14220 13596 14272
rect 16396 14220 16448 14272
rect 18052 14220 18104 14272
rect 18604 14220 18656 14272
rect 18972 14263 19024 14272
rect 18972 14229 18981 14263
rect 18981 14229 19015 14263
rect 19015 14229 19024 14263
rect 18972 14220 19024 14229
rect 22652 14560 22704 14612
rect 20444 14356 20496 14408
rect 19340 14288 19392 14340
rect 19800 14288 19852 14340
rect 20628 14220 20680 14272
rect 22100 14399 22152 14408
rect 22100 14365 22109 14399
rect 22109 14365 22143 14399
rect 22143 14365 22152 14399
rect 22100 14356 22152 14365
rect 22284 14356 22336 14408
rect 22560 14288 22612 14340
rect 23388 14288 23440 14340
rect 21180 14220 21232 14272
rect 2658 14118 2710 14170
rect 2722 14118 2774 14170
rect 2786 14118 2838 14170
rect 2850 14118 2902 14170
rect 2914 14118 2966 14170
rect 2978 14118 3030 14170
rect 8658 14118 8710 14170
rect 8722 14118 8774 14170
rect 8786 14118 8838 14170
rect 8850 14118 8902 14170
rect 8914 14118 8966 14170
rect 8978 14118 9030 14170
rect 14658 14118 14710 14170
rect 14722 14118 14774 14170
rect 14786 14118 14838 14170
rect 14850 14118 14902 14170
rect 14914 14118 14966 14170
rect 14978 14118 15030 14170
rect 20658 14118 20710 14170
rect 20722 14118 20774 14170
rect 20786 14118 20838 14170
rect 20850 14118 20902 14170
rect 20914 14118 20966 14170
rect 20978 14118 21030 14170
rect 6828 14016 6880 14068
rect 3700 13948 3752 14000
rect 1768 13880 1820 13932
rect 2136 13923 2188 13932
rect 2136 13889 2170 13923
rect 2170 13889 2188 13923
rect 2136 13880 2188 13889
rect 3148 13880 3200 13932
rect 3332 13923 3384 13932
rect 3332 13889 3341 13923
rect 3341 13889 3375 13923
rect 3375 13889 3384 13923
rect 3332 13880 3384 13889
rect 3884 13880 3936 13932
rect 4436 13880 4488 13932
rect 5080 13923 5132 13932
rect 5080 13889 5114 13923
rect 5114 13889 5132 13923
rect 5080 13880 5132 13889
rect 5632 13880 5684 13932
rect 4804 13855 4856 13864
rect 4804 13821 4813 13855
rect 4813 13821 4847 13855
rect 4847 13821 4856 13855
rect 4804 13812 4856 13821
rect 12992 14016 13044 14068
rect 13360 14016 13412 14068
rect 14188 14016 14240 14068
rect 16396 14016 16448 14068
rect 16488 14059 16540 14068
rect 16488 14025 16497 14059
rect 16497 14025 16531 14059
rect 16531 14025 16540 14059
rect 16488 14016 16540 14025
rect 9128 13880 9180 13932
rect 3056 13676 3108 13728
rect 6368 13744 6420 13796
rect 8392 13812 8444 13864
rect 9864 13948 9916 14000
rect 9956 13948 10008 14000
rect 11888 13948 11940 14000
rect 11980 13948 12032 14000
rect 11060 13923 11112 13932
rect 11060 13889 11078 13923
rect 11078 13889 11112 13923
rect 11060 13880 11112 13889
rect 11336 13855 11388 13864
rect 11336 13821 11345 13855
rect 11345 13821 11379 13855
rect 11379 13821 11388 13855
rect 11336 13812 11388 13821
rect 12900 13948 12952 14000
rect 13544 13991 13596 14000
rect 13544 13957 13553 13991
rect 13553 13957 13587 13991
rect 13587 13957 13596 13991
rect 13544 13948 13596 13957
rect 15108 13948 15160 14000
rect 12164 13880 12216 13932
rect 13820 13880 13872 13932
rect 17224 14016 17276 14068
rect 17684 14059 17736 14068
rect 17684 14025 17693 14059
rect 17693 14025 17727 14059
rect 17727 14025 17736 14059
rect 17684 14016 17736 14025
rect 18144 14016 18196 14068
rect 18236 14016 18288 14068
rect 19340 14016 19392 14068
rect 21272 14016 21324 14068
rect 22100 14016 22152 14068
rect 17040 13880 17092 13932
rect 18512 13948 18564 14000
rect 22652 13948 22704 14000
rect 23204 13948 23256 14000
rect 23296 13948 23348 14000
rect 11612 13744 11664 13796
rect 13820 13744 13872 13796
rect 17132 13744 17184 13796
rect 18052 13812 18104 13864
rect 19984 13880 20036 13932
rect 21456 13880 21508 13932
rect 21548 13923 21600 13932
rect 21548 13889 21557 13923
rect 21557 13889 21591 13923
rect 21591 13889 21600 13923
rect 21548 13880 21600 13889
rect 21732 13880 21784 13932
rect 21180 13812 21232 13864
rect 21364 13812 21416 13864
rect 14832 13719 14884 13728
rect 14832 13685 14841 13719
rect 14841 13685 14875 13719
rect 14875 13685 14884 13719
rect 14832 13676 14884 13685
rect 20812 13676 20864 13728
rect 1918 13574 1970 13626
rect 1982 13574 2034 13626
rect 2046 13574 2098 13626
rect 2110 13574 2162 13626
rect 2174 13574 2226 13626
rect 2238 13574 2290 13626
rect 7918 13574 7970 13626
rect 7982 13574 8034 13626
rect 8046 13574 8098 13626
rect 8110 13574 8162 13626
rect 8174 13574 8226 13626
rect 8238 13574 8290 13626
rect 13918 13574 13970 13626
rect 13982 13574 14034 13626
rect 14046 13574 14098 13626
rect 14110 13574 14162 13626
rect 14174 13574 14226 13626
rect 14238 13574 14290 13626
rect 19918 13574 19970 13626
rect 19982 13574 20034 13626
rect 20046 13574 20098 13626
rect 20110 13574 20162 13626
rect 20174 13574 20226 13626
rect 20238 13574 20290 13626
rect 3240 13472 3292 13524
rect 940 13336 992 13388
rect 3056 13268 3108 13320
rect 3516 13268 3568 13320
rect 7012 13404 7064 13456
rect 10784 13515 10836 13524
rect 10784 13481 10793 13515
rect 10793 13481 10827 13515
rect 10827 13481 10836 13515
rect 10784 13472 10836 13481
rect 12900 13472 12952 13524
rect 12992 13472 13044 13524
rect 9680 13404 9732 13456
rect 4068 13379 4120 13388
rect 4068 13345 4077 13379
rect 4077 13345 4111 13379
rect 4111 13345 4120 13379
rect 4068 13336 4120 13345
rect 13176 13379 13228 13388
rect 13176 13345 13185 13379
rect 13185 13345 13219 13379
rect 13219 13345 13228 13379
rect 13176 13336 13228 13345
rect 3240 13200 3292 13252
rect 3332 13243 3384 13252
rect 3332 13209 3350 13243
rect 3350 13209 3384 13243
rect 3332 13200 3384 13209
rect 4344 13243 4396 13252
rect 4344 13209 4378 13243
rect 4378 13209 4396 13243
rect 4344 13200 4396 13209
rect 6644 13268 6696 13320
rect 11152 13268 11204 13320
rect 11244 13268 11296 13320
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 11888 13268 11940 13320
rect 13452 13311 13504 13320
rect 13452 13277 13461 13311
rect 13461 13277 13495 13311
rect 13495 13277 13504 13311
rect 13452 13268 13504 13277
rect 14372 13472 14424 13524
rect 15384 13404 15436 13456
rect 15936 13472 15988 13524
rect 19892 13472 19944 13524
rect 22192 13472 22244 13524
rect 16396 13404 16448 13456
rect 14832 13336 14884 13388
rect 23388 13379 23440 13388
rect 23388 13345 23397 13379
rect 23397 13345 23431 13379
rect 23431 13345 23440 13379
rect 23388 13336 23440 13345
rect 3148 13132 3200 13184
rect 5356 13132 5408 13184
rect 5448 13175 5500 13184
rect 5448 13141 5457 13175
rect 5457 13141 5491 13175
rect 5491 13141 5500 13175
rect 5448 13132 5500 13141
rect 5816 13243 5868 13252
rect 5816 13209 5850 13243
rect 5850 13209 5868 13243
rect 5816 13200 5868 13209
rect 8392 13200 8444 13252
rect 7196 13132 7248 13184
rect 9036 13200 9088 13252
rect 9312 13132 9364 13184
rect 9496 13132 9548 13184
rect 11152 13132 11204 13184
rect 13820 13200 13872 13252
rect 17040 13268 17092 13320
rect 17316 13311 17368 13320
rect 17316 13277 17325 13311
rect 17325 13277 17359 13311
rect 17359 13277 17368 13311
rect 17316 13268 17368 13277
rect 15476 13243 15528 13252
rect 15476 13209 15485 13243
rect 15485 13209 15519 13243
rect 15519 13209 15528 13243
rect 15476 13200 15528 13209
rect 15292 13132 15344 13184
rect 18052 13268 18104 13320
rect 17960 13200 18012 13252
rect 19340 13268 19392 13320
rect 21548 13268 21600 13320
rect 21824 13268 21876 13320
rect 22376 13268 22428 13320
rect 20812 13200 20864 13252
rect 18144 13132 18196 13184
rect 18880 13175 18932 13184
rect 18880 13141 18889 13175
rect 18889 13141 18923 13175
rect 18923 13141 18932 13175
rect 18880 13132 18932 13141
rect 19248 13175 19300 13184
rect 19248 13141 19257 13175
rect 19257 13141 19291 13175
rect 19291 13141 19300 13175
rect 19248 13132 19300 13141
rect 19984 13132 20036 13184
rect 23388 13200 23440 13252
rect 2658 13030 2710 13082
rect 2722 13030 2774 13082
rect 2786 13030 2838 13082
rect 2850 13030 2902 13082
rect 2914 13030 2966 13082
rect 2978 13030 3030 13082
rect 8658 13030 8710 13082
rect 8722 13030 8774 13082
rect 8786 13030 8838 13082
rect 8850 13030 8902 13082
rect 8914 13030 8966 13082
rect 8978 13030 9030 13082
rect 14658 13030 14710 13082
rect 14722 13030 14774 13082
rect 14786 13030 14838 13082
rect 14850 13030 14902 13082
rect 14914 13030 14966 13082
rect 14978 13030 15030 13082
rect 20658 13030 20710 13082
rect 20722 13030 20774 13082
rect 20786 13030 20838 13082
rect 20850 13030 20902 13082
rect 20914 13030 20966 13082
rect 20978 13030 21030 13082
rect 4804 12928 4856 12980
rect 5356 12928 5408 12980
rect 3148 12860 3200 12912
rect 2964 12835 3016 12844
rect 4712 12860 4764 12912
rect 2964 12801 2993 12835
rect 2993 12801 3016 12835
rect 2964 12792 3016 12801
rect 3424 12792 3476 12844
rect 4896 12792 4948 12844
rect 11336 12928 11388 12980
rect 12808 12971 12860 12980
rect 1768 12588 1820 12640
rect 3516 12588 3568 12640
rect 6828 12835 6880 12844
rect 6828 12801 6837 12835
rect 6837 12801 6871 12835
rect 6871 12801 6880 12835
rect 6828 12792 6880 12801
rect 7196 12792 7248 12844
rect 7656 12835 7708 12844
rect 7656 12801 7665 12835
rect 7665 12801 7699 12835
rect 7699 12801 7708 12835
rect 7656 12792 7708 12801
rect 6736 12724 6788 12776
rect 8392 12792 8444 12844
rect 4620 12656 4672 12708
rect 7656 12656 7708 12708
rect 6184 12631 6236 12640
rect 6184 12597 6193 12631
rect 6193 12597 6227 12631
rect 6227 12597 6236 12631
rect 6184 12588 6236 12597
rect 7472 12588 7524 12640
rect 7564 12631 7616 12640
rect 7564 12597 7573 12631
rect 7573 12597 7607 12631
rect 7607 12597 7616 12631
rect 7564 12588 7616 12597
rect 9772 12656 9824 12708
rect 12808 12937 12817 12971
rect 12817 12937 12851 12971
rect 12851 12937 12860 12971
rect 12808 12928 12860 12937
rect 16856 12928 16908 12980
rect 17040 12928 17092 12980
rect 18880 12928 18932 12980
rect 19248 12928 19300 12980
rect 19800 12971 19852 12980
rect 19800 12937 19809 12971
rect 19809 12937 19843 12971
rect 19843 12937 19852 12971
rect 19800 12928 19852 12937
rect 11336 12835 11388 12844
rect 11336 12801 11345 12835
rect 11345 12801 11379 12835
rect 11379 12801 11388 12835
rect 11336 12792 11388 12801
rect 11520 12835 11572 12844
rect 11520 12801 11529 12835
rect 11529 12801 11563 12835
rect 11563 12801 11572 12835
rect 11520 12792 11572 12801
rect 15200 12860 15252 12912
rect 13636 12835 13688 12844
rect 13636 12801 13645 12835
rect 13645 12801 13679 12835
rect 13679 12801 13688 12835
rect 13636 12792 13688 12801
rect 13912 12835 13964 12844
rect 13912 12801 13921 12835
rect 13921 12801 13955 12835
rect 13955 12801 13964 12835
rect 13912 12792 13964 12801
rect 11612 12724 11664 12776
rect 9404 12588 9456 12640
rect 11428 12656 11480 12708
rect 14280 12699 14332 12708
rect 14280 12665 14289 12699
rect 14289 12665 14323 12699
rect 14323 12665 14332 12699
rect 14280 12656 14332 12665
rect 15108 12792 15160 12844
rect 16672 12724 16724 12776
rect 16212 12699 16264 12708
rect 16212 12665 16221 12699
rect 16221 12665 16255 12699
rect 16255 12665 16264 12699
rect 16212 12656 16264 12665
rect 16948 12792 17000 12844
rect 19616 12792 19668 12844
rect 21640 12860 21692 12912
rect 22192 12860 22244 12912
rect 19892 12792 19944 12844
rect 21088 12792 21140 12844
rect 21364 12792 21416 12844
rect 22376 12792 22428 12844
rect 19984 12724 20036 12776
rect 21732 12724 21784 12776
rect 16856 12656 16908 12708
rect 11152 12631 11204 12640
rect 11152 12597 11161 12631
rect 11161 12597 11195 12631
rect 11195 12597 11204 12631
rect 11152 12588 11204 12597
rect 11336 12588 11388 12640
rect 11796 12588 11848 12640
rect 13728 12588 13780 12640
rect 14372 12631 14424 12640
rect 14372 12597 14381 12631
rect 14381 12597 14415 12631
rect 14415 12597 14424 12631
rect 14372 12588 14424 12597
rect 17592 12588 17644 12640
rect 20444 12588 20496 12640
rect 21732 12588 21784 12640
rect 22836 12724 22888 12776
rect 22560 12588 22612 12640
rect 1918 12486 1970 12538
rect 1982 12486 2034 12538
rect 2046 12486 2098 12538
rect 2110 12486 2162 12538
rect 2174 12486 2226 12538
rect 2238 12486 2290 12538
rect 7918 12486 7970 12538
rect 7982 12486 8034 12538
rect 8046 12486 8098 12538
rect 8110 12486 8162 12538
rect 8174 12486 8226 12538
rect 8238 12486 8290 12538
rect 13918 12486 13970 12538
rect 13982 12486 14034 12538
rect 14046 12486 14098 12538
rect 14110 12486 14162 12538
rect 14174 12486 14226 12538
rect 14238 12486 14290 12538
rect 19918 12486 19970 12538
rect 19982 12486 20034 12538
rect 20046 12486 20098 12538
rect 20110 12486 20162 12538
rect 20174 12486 20226 12538
rect 20238 12486 20290 12538
rect 3332 12384 3384 12436
rect 7656 12384 7708 12436
rect 10232 12384 10284 12436
rect 13452 12384 13504 12436
rect 13544 12384 13596 12436
rect 14556 12384 14608 12436
rect 15292 12384 15344 12436
rect 12348 12316 12400 12368
rect 1400 12248 1452 12300
rect 4344 12291 4396 12300
rect 4344 12257 4353 12291
rect 4353 12257 4387 12291
rect 4387 12257 4396 12291
rect 4344 12248 4396 12257
rect 9404 12248 9456 12300
rect 13452 12291 13504 12300
rect 13452 12257 13461 12291
rect 13461 12257 13495 12291
rect 13495 12257 13504 12291
rect 13452 12248 13504 12257
rect 940 12180 992 12232
rect 3332 12180 3384 12232
rect 3976 12112 4028 12164
rect 4160 12112 4212 12164
rect 4896 12112 4948 12164
rect 7196 12112 7248 12164
rect 8392 12112 8444 12164
rect 8944 12223 8996 12232
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 9864 12180 9916 12232
rect 9220 12112 9272 12164
rect 13360 12180 13412 12232
rect 18144 12316 18196 12368
rect 6276 12044 6328 12096
rect 7472 12044 7524 12096
rect 11888 12112 11940 12164
rect 17500 12248 17552 12300
rect 17592 12248 17644 12300
rect 10232 12087 10284 12096
rect 10232 12053 10241 12087
rect 10241 12053 10275 12087
rect 10275 12053 10284 12087
rect 10232 12044 10284 12053
rect 11336 12044 11388 12096
rect 13636 12044 13688 12096
rect 14372 12044 14424 12096
rect 16028 12223 16080 12232
rect 16028 12189 16037 12223
rect 16037 12189 16071 12223
rect 16071 12189 16080 12223
rect 16028 12180 16080 12189
rect 18144 12180 18196 12232
rect 16672 12112 16724 12164
rect 19064 12223 19116 12232
rect 19064 12189 19073 12223
rect 19073 12189 19107 12223
rect 19107 12189 19116 12223
rect 19064 12180 19116 12189
rect 23112 12384 23164 12436
rect 23388 12384 23440 12436
rect 21180 12248 21232 12300
rect 21824 12248 21876 12300
rect 19708 12180 19760 12232
rect 23480 12180 23532 12232
rect 16120 12044 16172 12096
rect 18420 12044 18472 12096
rect 20444 12112 20496 12164
rect 20536 12087 20588 12096
rect 20536 12053 20545 12087
rect 20545 12053 20579 12087
rect 20579 12053 20588 12087
rect 20536 12044 20588 12053
rect 21088 12044 21140 12096
rect 22836 12044 22888 12096
rect 2658 11942 2710 11994
rect 2722 11942 2774 11994
rect 2786 11942 2838 11994
rect 2850 11942 2902 11994
rect 2914 11942 2966 11994
rect 2978 11942 3030 11994
rect 8658 11942 8710 11994
rect 8722 11942 8774 11994
rect 8786 11942 8838 11994
rect 8850 11942 8902 11994
rect 8914 11942 8966 11994
rect 8978 11942 9030 11994
rect 14658 11942 14710 11994
rect 14722 11942 14774 11994
rect 14786 11942 14838 11994
rect 14850 11942 14902 11994
rect 14914 11942 14966 11994
rect 14978 11942 15030 11994
rect 20658 11942 20710 11994
rect 20722 11942 20774 11994
rect 20786 11942 20838 11994
rect 20850 11942 20902 11994
rect 20914 11942 20966 11994
rect 20978 11942 21030 11994
rect 1584 11840 1636 11892
rect 11060 11840 11112 11892
rect 1768 11772 1820 11824
rect 2504 11772 2556 11824
rect 9772 11772 9824 11824
rect 3240 11704 3292 11756
rect 5908 11747 5960 11756
rect 5908 11713 5937 11747
rect 5937 11713 5960 11747
rect 5908 11704 5960 11713
rect 6092 11704 6144 11756
rect 1492 11636 1544 11688
rect 3056 11636 3108 11688
rect 6368 11679 6420 11688
rect 6368 11645 6377 11679
rect 6377 11645 6411 11679
rect 6411 11645 6420 11679
rect 6368 11636 6420 11645
rect 9680 11747 9732 11756
rect 9680 11713 9689 11747
rect 9689 11713 9723 11747
rect 9723 11713 9732 11747
rect 9680 11704 9732 11713
rect 10508 11704 10560 11756
rect 15752 11840 15804 11892
rect 12808 11772 12860 11824
rect 15108 11772 15160 11824
rect 11612 11747 11664 11756
rect 11612 11713 11621 11747
rect 11621 11713 11655 11747
rect 11655 11713 11664 11747
rect 11612 11704 11664 11713
rect 11704 11704 11756 11756
rect 15568 11704 15620 11756
rect 21088 11840 21140 11892
rect 21548 11883 21600 11892
rect 21548 11849 21557 11883
rect 21557 11849 21591 11883
rect 21591 11849 21600 11883
rect 21548 11840 21600 11849
rect 21640 11840 21692 11892
rect 20536 11772 20588 11824
rect 21364 11772 21416 11824
rect 22560 11772 22612 11824
rect 18604 11704 18656 11756
rect 1768 11611 1820 11620
rect 1768 11577 1777 11611
rect 1777 11577 1811 11611
rect 1811 11577 1820 11611
rect 1768 11568 1820 11577
rect 4344 11568 4396 11620
rect 11244 11636 11296 11688
rect 21640 11747 21692 11756
rect 21640 11713 21649 11747
rect 21649 11713 21683 11747
rect 21683 11713 21692 11747
rect 21640 11704 21692 11713
rect 21916 11704 21968 11756
rect 23296 11747 23348 11756
rect 23296 11713 23305 11747
rect 23305 11713 23339 11747
rect 23339 11713 23348 11747
rect 23296 11704 23348 11713
rect 3332 11500 3384 11552
rect 3516 11500 3568 11552
rect 7656 11500 7708 11552
rect 8484 11500 8536 11552
rect 9128 11543 9180 11552
rect 9128 11509 9137 11543
rect 9137 11509 9171 11543
rect 9171 11509 9180 11543
rect 9128 11500 9180 11509
rect 11152 11500 11204 11552
rect 11796 11500 11848 11552
rect 12992 11543 13044 11552
rect 12992 11509 13001 11543
rect 13001 11509 13035 11543
rect 13035 11509 13044 11543
rect 12992 11500 13044 11509
rect 17592 11568 17644 11620
rect 16212 11500 16264 11552
rect 16764 11500 16816 11552
rect 19800 11500 19852 11552
rect 21180 11500 21232 11552
rect 21824 11679 21876 11688
rect 21824 11645 21833 11679
rect 21833 11645 21867 11679
rect 21867 11645 21876 11679
rect 21824 11636 21876 11645
rect 23020 11568 23072 11620
rect 22468 11500 22520 11552
rect 1918 11398 1970 11450
rect 1982 11398 2034 11450
rect 2046 11398 2098 11450
rect 2110 11398 2162 11450
rect 2174 11398 2226 11450
rect 2238 11398 2290 11450
rect 7918 11398 7970 11450
rect 7982 11398 8034 11450
rect 8046 11398 8098 11450
rect 8110 11398 8162 11450
rect 8174 11398 8226 11450
rect 8238 11398 8290 11450
rect 13918 11398 13970 11450
rect 13982 11398 14034 11450
rect 14046 11398 14098 11450
rect 14110 11398 14162 11450
rect 14174 11398 14226 11450
rect 14238 11398 14290 11450
rect 19918 11398 19970 11450
rect 19982 11398 20034 11450
rect 20046 11398 20098 11450
rect 20110 11398 20162 11450
rect 20174 11398 20226 11450
rect 20238 11398 20290 11450
rect 5632 11296 5684 11348
rect 11704 11296 11756 11348
rect 12808 11296 12860 11348
rect 13268 11296 13320 11348
rect 11612 11228 11664 11280
rect 15476 11296 15528 11348
rect 3332 11160 3384 11212
rect 3608 11160 3660 11212
rect 2320 11092 2372 11144
rect 4436 11135 4488 11144
rect 4436 11101 4445 11135
rect 4445 11101 4479 11135
rect 4479 11101 4488 11135
rect 4436 11092 4488 11101
rect 5816 11160 5868 11212
rect 14096 11160 14148 11212
rect 15292 11271 15344 11280
rect 15292 11237 15301 11271
rect 15301 11237 15335 11271
rect 15335 11237 15344 11271
rect 23296 11296 23348 11348
rect 15292 11228 15344 11237
rect 16672 11160 16724 11212
rect 17132 11203 17184 11212
rect 17132 11169 17141 11203
rect 17141 11169 17175 11203
rect 17175 11169 17184 11203
rect 17132 11160 17184 11169
rect 18512 11160 18564 11212
rect 19708 11203 19760 11212
rect 19708 11169 19717 11203
rect 19717 11169 19751 11203
rect 19751 11169 19760 11203
rect 19708 11160 19760 11169
rect 5448 11092 5500 11144
rect 5540 11092 5592 11144
rect 7380 11135 7432 11144
rect 7380 11101 7389 11135
rect 7389 11101 7423 11135
rect 7423 11101 7432 11135
rect 7380 11092 7432 11101
rect 7656 11135 7708 11144
rect 7656 11101 7690 11135
rect 7690 11101 7708 11135
rect 7656 11092 7708 11101
rect 10784 11092 10836 11144
rect 12992 11092 13044 11144
rect 13268 11135 13320 11144
rect 13268 11101 13286 11135
rect 13286 11101 13320 11135
rect 13268 11092 13320 11101
rect 13636 11135 13688 11144
rect 13636 11101 13645 11135
rect 13645 11101 13679 11135
rect 13679 11101 13688 11135
rect 13636 11092 13688 11101
rect 3240 11024 3292 11076
rect 3700 11024 3752 11076
rect 4528 11024 4580 11076
rect 4804 11024 4856 11076
rect 9128 11024 9180 11076
rect 9220 11024 9272 11076
rect 11152 11024 11204 11076
rect 7472 10956 7524 11008
rect 15108 11092 15160 11144
rect 14280 11024 14332 11076
rect 15384 11024 15436 11076
rect 16948 10956 17000 11008
rect 22008 11228 22060 11280
rect 21548 11203 21600 11212
rect 21548 11169 21557 11203
rect 21557 11169 21591 11203
rect 21591 11169 21600 11203
rect 21548 11160 21600 11169
rect 20352 11092 20404 11144
rect 22100 11024 22152 11076
rect 17776 10956 17828 11008
rect 19616 10956 19668 11008
rect 21456 10956 21508 11008
rect 22008 10956 22060 11008
rect 23020 11135 23072 11144
rect 23020 11101 23029 11135
rect 23029 11101 23063 11135
rect 23063 11101 23072 11135
rect 23020 11092 23072 11101
rect 23112 11135 23164 11144
rect 23112 11101 23121 11135
rect 23121 11101 23155 11135
rect 23155 11101 23164 11135
rect 23112 11092 23164 11101
rect 2658 10854 2710 10906
rect 2722 10854 2774 10906
rect 2786 10854 2838 10906
rect 2850 10854 2902 10906
rect 2914 10854 2966 10906
rect 2978 10854 3030 10906
rect 8658 10854 8710 10906
rect 8722 10854 8774 10906
rect 8786 10854 8838 10906
rect 8850 10854 8902 10906
rect 8914 10854 8966 10906
rect 8978 10854 9030 10906
rect 14658 10854 14710 10906
rect 14722 10854 14774 10906
rect 14786 10854 14838 10906
rect 14850 10854 14902 10906
rect 14914 10854 14966 10906
rect 14978 10854 15030 10906
rect 20658 10854 20710 10906
rect 20722 10854 20774 10906
rect 20786 10854 20838 10906
rect 20850 10854 20902 10906
rect 20914 10854 20966 10906
rect 20978 10854 21030 10906
rect 1216 10616 1268 10668
rect 2228 10684 2280 10736
rect 2504 10684 2556 10736
rect 5540 10752 5592 10804
rect 1860 10616 1912 10668
rect 2596 10616 2648 10668
rect 3148 10616 3200 10668
rect 3332 10616 3384 10668
rect 7288 10684 7340 10736
rect 7472 10684 7524 10736
rect 8484 10727 8536 10736
rect 8484 10693 8493 10727
rect 8493 10693 8527 10727
rect 8527 10693 8536 10727
rect 8484 10684 8536 10693
rect 3884 10616 3936 10668
rect 6460 10659 6512 10668
rect 6460 10625 6469 10659
rect 6469 10625 6503 10659
rect 6503 10625 6512 10659
rect 6460 10616 6512 10625
rect 7840 10616 7892 10668
rect 13820 10752 13872 10804
rect 15568 10752 15620 10804
rect 16580 10752 16632 10804
rect 17316 10752 17368 10804
rect 17500 10752 17552 10804
rect 4252 10548 4304 10600
rect 16672 10684 16724 10736
rect 11612 10659 11664 10668
rect 11612 10625 11621 10659
rect 11621 10625 11655 10659
rect 11655 10625 11664 10659
rect 11612 10616 11664 10625
rect 13636 10616 13688 10668
rect 13728 10659 13780 10668
rect 13728 10625 13737 10659
rect 13737 10625 13771 10659
rect 13771 10625 13780 10659
rect 13728 10616 13780 10625
rect 13820 10616 13872 10668
rect 14372 10659 14424 10668
rect 14372 10625 14406 10659
rect 14406 10625 14424 10659
rect 14372 10616 14424 10625
rect 14648 10616 14700 10668
rect 16120 10616 16172 10668
rect 17960 10684 18012 10736
rect 18420 10684 18472 10736
rect 18972 10684 19024 10736
rect 11520 10480 11572 10532
rect 14096 10591 14148 10600
rect 14096 10557 14105 10591
rect 14105 10557 14139 10591
rect 14139 10557 14148 10591
rect 14096 10548 14148 10557
rect 16580 10548 16632 10600
rect 19432 10616 19484 10668
rect 17224 10548 17276 10600
rect 5080 10412 5132 10464
rect 6920 10412 6972 10464
rect 10324 10412 10376 10464
rect 10416 10455 10468 10464
rect 10416 10421 10425 10455
rect 10425 10421 10459 10455
rect 10459 10421 10468 10455
rect 10416 10412 10468 10421
rect 12532 10412 12584 10464
rect 19064 10480 19116 10532
rect 20444 10616 20496 10668
rect 21364 10659 21416 10668
rect 21364 10625 21373 10659
rect 21373 10625 21407 10659
rect 21407 10625 21416 10659
rect 21364 10616 21416 10625
rect 21916 10616 21968 10668
rect 22376 10752 22428 10804
rect 22928 10752 22980 10804
rect 23020 10752 23072 10804
rect 23204 10659 23256 10668
rect 23204 10625 23213 10659
rect 23213 10625 23247 10659
rect 23247 10625 23256 10659
rect 23204 10616 23256 10625
rect 20904 10548 20956 10600
rect 14464 10412 14516 10464
rect 19156 10412 19208 10464
rect 21640 10548 21692 10600
rect 1918 10310 1970 10362
rect 1982 10310 2034 10362
rect 2046 10310 2098 10362
rect 2110 10310 2162 10362
rect 2174 10310 2226 10362
rect 2238 10310 2290 10362
rect 7918 10310 7970 10362
rect 7982 10310 8034 10362
rect 8046 10310 8098 10362
rect 8110 10310 8162 10362
rect 8174 10310 8226 10362
rect 8238 10310 8290 10362
rect 13918 10310 13970 10362
rect 13982 10310 14034 10362
rect 14046 10310 14098 10362
rect 14110 10310 14162 10362
rect 14174 10310 14226 10362
rect 14238 10310 14290 10362
rect 19918 10310 19970 10362
rect 19982 10310 20034 10362
rect 20046 10310 20098 10362
rect 20110 10310 20162 10362
rect 20174 10310 20226 10362
rect 20238 10310 20290 10362
rect 1584 10208 1636 10260
rect 2504 10208 2556 10260
rect 3516 10140 3568 10192
rect 3884 10140 3936 10192
rect 6368 10208 6420 10260
rect 7196 10208 7248 10260
rect 7748 10140 7800 10192
rect 2228 10004 2280 10056
rect 2596 10004 2648 10056
rect 1308 9868 1360 9920
rect 4344 10072 4396 10124
rect 7840 10072 7892 10124
rect 10600 10140 10652 10192
rect 13636 10208 13688 10260
rect 17776 10208 17828 10260
rect 9864 10072 9916 10124
rect 11152 10072 11204 10124
rect 4528 9936 4580 9988
rect 5540 9936 5592 9988
rect 6000 9936 6052 9988
rect 4712 9868 4764 9920
rect 9312 9936 9364 9988
rect 11520 10004 11572 10056
rect 11796 10004 11848 10056
rect 14188 10072 14240 10124
rect 20352 10208 20404 10260
rect 18880 10140 18932 10192
rect 12532 10047 12584 10056
rect 12532 10013 12541 10047
rect 12541 10013 12575 10047
rect 12575 10013 12584 10047
rect 12532 10004 12584 10013
rect 12808 10047 12860 10056
rect 12808 10013 12842 10047
rect 12842 10013 12860 10047
rect 12808 10004 12860 10013
rect 15568 10047 15620 10056
rect 15568 10013 15577 10047
rect 15577 10013 15611 10047
rect 15611 10013 15620 10047
rect 15568 10004 15620 10013
rect 19340 10004 19392 10056
rect 20076 10004 20128 10056
rect 21456 10004 21508 10056
rect 23296 10115 23348 10124
rect 23296 10081 23305 10115
rect 23305 10081 23339 10115
rect 23339 10081 23348 10115
rect 23296 10072 23348 10081
rect 22008 10004 22060 10056
rect 12624 9936 12676 9988
rect 14096 9936 14148 9988
rect 17592 9936 17644 9988
rect 18144 9936 18196 9988
rect 18236 9979 18288 9988
rect 18236 9945 18254 9979
rect 18254 9945 18288 9979
rect 18236 9936 18288 9945
rect 18512 9936 18564 9988
rect 19156 9936 19208 9988
rect 21916 9936 21968 9988
rect 6276 9868 6328 9920
rect 8484 9868 8536 9920
rect 10692 9868 10744 9920
rect 11612 9868 11664 9920
rect 12532 9868 12584 9920
rect 17132 9911 17184 9920
rect 17132 9877 17141 9911
rect 17141 9877 17175 9911
rect 17175 9877 17184 9911
rect 17132 9868 17184 9877
rect 20904 9868 20956 9920
rect 21640 9868 21692 9920
rect 22468 10047 22520 10056
rect 22468 10013 22477 10047
rect 22477 10013 22511 10047
rect 22511 10013 22520 10047
rect 22468 10004 22520 10013
rect 22744 10004 22796 10056
rect 2658 9766 2710 9818
rect 2722 9766 2774 9818
rect 2786 9766 2838 9818
rect 2850 9766 2902 9818
rect 2914 9766 2966 9818
rect 2978 9766 3030 9818
rect 8658 9766 8710 9818
rect 8722 9766 8774 9818
rect 8786 9766 8838 9818
rect 8850 9766 8902 9818
rect 8914 9766 8966 9818
rect 8978 9766 9030 9818
rect 14658 9766 14710 9818
rect 14722 9766 14774 9818
rect 14786 9766 14838 9818
rect 14850 9766 14902 9818
rect 14914 9766 14966 9818
rect 14978 9766 15030 9818
rect 20658 9766 20710 9818
rect 20722 9766 20774 9818
rect 20786 9766 20838 9818
rect 20850 9766 20902 9818
rect 20914 9766 20966 9818
rect 20978 9766 21030 9818
rect 2228 9664 2280 9716
rect 6000 9664 6052 9716
rect 6736 9664 6788 9716
rect 10324 9664 10376 9716
rect 14372 9664 14424 9716
rect 14464 9664 14516 9716
rect 21364 9664 21416 9716
rect 3332 9596 3384 9648
rect 6828 9596 6880 9648
rect 11980 9596 12032 9648
rect 14280 9596 14332 9648
rect 14648 9639 14700 9648
rect 14648 9605 14657 9639
rect 14657 9605 14691 9639
rect 14691 9605 14700 9639
rect 14648 9596 14700 9605
rect 15476 9596 15528 9648
rect 16396 9639 16448 9648
rect 16396 9605 16405 9639
rect 16405 9605 16439 9639
rect 16439 9605 16448 9639
rect 16396 9596 16448 9605
rect 16672 9639 16724 9648
rect 16672 9605 16681 9639
rect 16681 9605 16715 9639
rect 16715 9605 16724 9639
rect 16672 9596 16724 9605
rect 19524 9596 19576 9648
rect 2228 9571 2280 9580
rect 2228 9537 2237 9571
rect 2237 9537 2271 9571
rect 2271 9537 2280 9571
rect 2228 9528 2280 9537
rect 2964 9460 3016 9512
rect 4160 9528 4212 9580
rect 4620 9528 4672 9580
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 5080 9571 5132 9580
rect 5080 9537 5103 9571
rect 5103 9537 5132 9571
rect 5080 9528 5132 9537
rect 5540 9528 5592 9580
rect 3608 9460 3660 9512
rect 4804 9503 4856 9512
rect 4804 9469 4813 9503
rect 4813 9469 4847 9503
rect 4847 9469 4856 9503
rect 4804 9460 4856 9469
rect 2412 9435 2464 9444
rect 2412 9401 2421 9435
rect 2421 9401 2455 9435
rect 2455 9401 2464 9435
rect 2412 9392 2464 9401
rect 2596 9392 2648 9444
rect 3240 9324 3292 9376
rect 7104 9392 7156 9444
rect 7196 9324 7248 9376
rect 10416 9528 10468 9580
rect 9312 9460 9364 9512
rect 10600 9571 10652 9580
rect 10600 9537 10609 9571
rect 10609 9537 10643 9571
rect 10643 9537 10652 9571
rect 10600 9528 10652 9537
rect 11520 9528 11572 9580
rect 13452 9528 13504 9580
rect 14096 9528 14148 9580
rect 11704 9460 11756 9512
rect 12532 9503 12584 9512
rect 12532 9469 12541 9503
rect 12541 9469 12575 9503
rect 12575 9469 12584 9503
rect 12532 9460 12584 9469
rect 9312 9324 9364 9376
rect 12992 9392 13044 9444
rect 17868 9392 17920 9444
rect 9680 9324 9732 9376
rect 11244 9324 11296 9376
rect 11888 9324 11940 9376
rect 12808 9367 12860 9376
rect 12808 9333 12817 9367
rect 12817 9333 12851 9367
rect 12851 9333 12860 9367
rect 12808 9324 12860 9333
rect 14188 9324 14240 9376
rect 15384 9324 15436 9376
rect 17408 9324 17460 9376
rect 17960 9367 18012 9376
rect 17960 9333 17969 9367
rect 17969 9333 18003 9367
rect 18003 9333 18012 9367
rect 17960 9324 18012 9333
rect 20812 9528 20864 9580
rect 21916 9528 21968 9580
rect 23480 9571 23532 9580
rect 23480 9537 23489 9571
rect 23489 9537 23523 9571
rect 23523 9537 23532 9571
rect 23480 9528 23532 9537
rect 21364 9503 21416 9512
rect 21364 9469 21366 9503
rect 21366 9469 21400 9503
rect 21400 9469 21416 9503
rect 21364 9460 21416 9469
rect 21732 9460 21784 9512
rect 20352 9392 20404 9444
rect 23296 9435 23348 9444
rect 23296 9401 23305 9435
rect 23305 9401 23339 9435
rect 23339 9401 23348 9435
rect 23296 9392 23348 9401
rect 23112 9324 23164 9376
rect 1918 9222 1970 9274
rect 1982 9222 2034 9274
rect 2046 9222 2098 9274
rect 2110 9222 2162 9274
rect 2174 9222 2226 9274
rect 2238 9222 2290 9274
rect 7918 9222 7970 9274
rect 7982 9222 8034 9274
rect 8046 9222 8098 9274
rect 8110 9222 8162 9274
rect 8174 9222 8226 9274
rect 8238 9222 8290 9274
rect 13918 9222 13970 9274
rect 13982 9222 14034 9274
rect 14046 9222 14098 9274
rect 14110 9222 14162 9274
rect 14174 9222 14226 9274
rect 14238 9222 14290 9274
rect 19918 9222 19970 9274
rect 19982 9222 20034 9274
rect 20046 9222 20098 9274
rect 20110 9222 20162 9274
rect 20174 9222 20226 9274
rect 20238 9222 20290 9274
rect 5080 9120 5132 9172
rect 8392 9120 8444 9172
rect 9864 9120 9916 9172
rect 11980 9163 12032 9172
rect 11980 9129 11989 9163
rect 11989 9129 12023 9163
rect 12023 9129 12032 9163
rect 11980 9120 12032 9129
rect 12532 9163 12584 9172
rect 12532 9129 12541 9163
rect 12541 9129 12575 9163
rect 12575 9129 12584 9163
rect 12532 9120 12584 9129
rect 12808 9120 12860 9172
rect 2136 8916 2188 8968
rect 1860 8848 1912 8900
rect 2964 8916 3016 8968
rect 3516 8916 3568 8968
rect 3976 8916 4028 8968
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 4712 8916 4764 8968
rect 5080 8916 5132 8968
rect 8484 8916 8536 8968
rect 9220 9052 9272 9104
rect 17408 9163 17460 9172
rect 17408 9129 17417 9163
rect 17417 9129 17451 9163
rect 17451 9129 17460 9163
rect 17408 9120 17460 9129
rect 19156 9120 19208 9172
rect 17592 8984 17644 9036
rect 18604 9052 18656 9104
rect 19248 9052 19300 9104
rect 20352 9052 20404 9104
rect 20536 9052 20588 9104
rect 4344 8891 4396 8900
rect 4344 8857 4378 8891
rect 4378 8857 4396 8891
rect 4344 8848 4396 8857
rect 3608 8823 3660 8832
rect 3608 8789 3617 8823
rect 3617 8789 3651 8823
rect 3651 8789 3660 8823
rect 3608 8780 3660 8789
rect 5632 8848 5684 8900
rect 5448 8823 5500 8832
rect 5448 8789 5457 8823
rect 5457 8789 5491 8823
rect 5491 8789 5500 8823
rect 5448 8780 5500 8789
rect 6552 8780 6604 8832
rect 8576 8848 8628 8900
rect 9220 8959 9272 8968
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 9312 8916 9364 8968
rect 13820 8916 13872 8968
rect 13912 8959 13964 8968
rect 13912 8925 13921 8959
rect 13921 8925 13955 8959
rect 13955 8925 13964 8959
rect 13912 8916 13964 8925
rect 14188 8916 14240 8968
rect 9864 8848 9916 8900
rect 13544 8848 13596 8900
rect 14556 8848 14608 8900
rect 17960 8848 18012 8900
rect 10232 8780 10284 8832
rect 13820 8780 13872 8832
rect 14648 8780 14700 8832
rect 18512 8891 18564 8900
rect 18512 8857 18521 8891
rect 18521 8857 18555 8891
rect 18555 8857 18564 8891
rect 18512 8848 18564 8857
rect 18696 8848 18748 8900
rect 18788 8780 18840 8832
rect 22652 8984 22704 9036
rect 21364 8916 21416 8968
rect 22100 8823 22152 8832
rect 22100 8789 22109 8823
rect 22109 8789 22143 8823
rect 22143 8789 22152 8823
rect 22100 8780 22152 8789
rect 23296 8780 23348 8832
rect 2658 8678 2710 8730
rect 2722 8678 2774 8730
rect 2786 8678 2838 8730
rect 2850 8678 2902 8730
rect 2914 8678 2966 8730
rect 2978 8678 3030 8730
rect 8658 8678 8710 8730
rect 8722 8678 8774 8730
rect 8786 8678 8838 8730
rect 8850 8678 8902 8730
rect 8914 8678 8966 8730
rect 8978 8678 9030 8730
rect 14658 8678 14710 8730
rect 14722 8678 14774 8730
rect 14786 8678 14838 8730
rect 14850 8678 14902 8730
rect 14914 8678 14966 8730
rect 14978 8678 15030 8730
rect 20658 8678 20710 8730
rect 20722 8678 20774 8730
rect 20786 8678 20838 8730
rect 20850 8678 20902 8730
rect 20914 8678 20966 8730
rect 20978 8678 21030 8730
rect 9220 8576 9272 8628
rect 13912 8576 13964 8628
rect 2504 8508 2556 8560
rect 3332 8508 3384 8560
rect 3608 8551 3660 8560
rect 3608 8517 3642 8551
rect 3642 8517 3660 8551
rect 3608 8508 3660 8517
rect 3700 8508 3752 8560
rect 3976 8508 4028 8560
rect 5172 8508 5224 8560
rect 7196 8508 7248 8560
rect 7840 8508 7892 8560
rect 9680 8508 9732 8560
rect 14188 8551 14240 8560
rect 14188 8517 14197 8551
rect 14197 8517 14231 8551
rect 14231 8517 14240 8551
rect 14188 8508 14240 8517
rect 1860 8440 1912 8492
rect 2136 8440 2188 8492
rect 5540 8440 5592 8492
rect 3240 8415 3292 8424
rect 3240 8381 3249 8415
rect 3249 8381 3283 8415
rect 3283 8381 3292 8415
rect 3240 8372 3292 8381
rect 3332 8415 3384 8424
rect 3332 8381 3341 8415
rect 3341 8381 3375 8415
rect 3375 8381 3384 8415
rect 3332 8372 3384 8381
rect 6184 8415 6236 8424
rect 6184 8381 6193 8415
rect 6193 8381 6227 8415
rect 6227 8381 6236 8415
rect 6184 8372 6236 8381
rect 12440 8483 12492 8492
rect 12440 8449 12449 8483
rect 12449 8449 12483 8483
rect 12483 8449 12492 8483
rect 12440 8440 12492 8449
rect 15292 8576 15344 8628
rect 16120 8576 16172 8628
rect 16212 8619 16264 8628
rect 16212 8585 16221 8619
rect 16221 8585 16255 8619
rect 16255 8585 16264 8619
rect 16212 8576 16264 8585
rect 19064 8576 19116 8628
rect 21272 8576 21324 8628
rect 21824 8576 21876 8628
rect 22192 8576 22244 8628
rect 18512 8508 18564 8560
rect 20536 8508 20588 8560
rect 15384 8440 15436 8492
rect 15752 8483 15804 8492
rect 15752 8449 15770 8483
rect 15770 8449 15804 8483
rect 15752 8440 15804 8449
rect 16304 8483 16356 8492
rect 16304 8449 16313 8483
rect 16313 8449 16347 8483
rect 16347 8449 16356 8483
rect 16304 8440 16356 8449
rect 17132 8440 17184 8492
rect 8944 8372 8996 8424
rect 13728 8372 13780 8424
rect 3516 8236 3568 8288
rect 3608 8236 3660 8288
rect 4528 8236 4580 8288
rect 4896 8236 4948 8288
rect 15016 8372 15068 8424
rect 16580 8372 16632 8424
rect 17960 8483 18012 8492
rect 17960 8449 17969 8483
rect 17969 8449 18003 8483
rect 18003 8449 18012 8483
rect 17960 8440 18012 8449
rect 18880 8372 18932 8424
rect 19800 8372 19852 8424
rect 5908 8236 5960 8288
rect 6460 8236 6512 8288
rect 10048 8279 10100 8288
rect 10048 8245 10057 8279
rect 10057 8245 10091 8279
rect 10091 8245 10100 8279
rect 10048 8236 10100 8245
rect 16120 8304 16172 8356
rect 16672 8304 16724 8356
rect 16396 8236 16448 8288
rect 18236 8304 18288 8356
rect 20444 8440 20496 8492
rect 21640 8440 21692 8492
rect 21732 8440 21784 8492
rect 23296 8483 23348 8492
rect 23296 8449 23305 8483
rect 23305 8449 23339 8483
rect 23339 8449 23348 8483
rect 23296 8440 23348 8449
rect 21180 8236 21232 8288
rect 22468 8236 22520 8288
rect 1918 8134 1970 8186
rect 1982 8134 2034 8186
rect 2046 8134 2098 8186
rect 2110 8134 2162 8186
rect 2174 8134 2226 8186
rect 2238 8134 2290 8186
rect 7918 8134 7970 8186
rect 7982 8134 8034 8186
rect 8046 8134 8098 8186
rect 8110 8134 8162 8186
rect 8174 8134 8226 8186
rect 8238 8134 8290 8186
rect 13918 8134 13970 8186
rect 13982 8134 14034 8186
rect 14046 8134 14098 8186
rect 14110 8134 14162 8186
rect 14174 8134 14226 8186
rect 14238 8134 14290 8186
rect 19918 8134 19970 8186
rect 19982 8134 20034 8186
rect 20046 8134 20098 8186
rect 20110 8134 20162 8186
rect 20174 8134 20226 8186
rect 20238 8134 20290 8186
rect 2228 8032 2280 8084
rect 2412 8032 2464 8084
rect 3516 8032 3568 8084
rect 3608 8075 3660 8084
rect 3608 8041 3617 8075
rect 3617 8041 3651 8075
rect 3651 8041 3660 8075
rect 3608 8032 3660 8041
rect 5172 8032 5224 8084
rect 8944 8075 8996 8084
rect 8944 8041 8953 8075
rect 8953 8041 8987 8075
rect 8987 8041 8996 8075
rect 8944 8032 8996 8041
rect 9404 8032 9456 8084
rect 14280 8032 14332 8084
rect 14464 8032 14516 8084
rect 16396 8032 16448 8084
rect 10508 7964 10560 8016
rect 11980 7964 12032 8016
rect 10692 7939 10744 7948
rect 2320 7828 2372 7880
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 4896 7828 4948 7880
rect 5448 7871 5500 7880
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 2596 7760 2648 7812
rect 3148 7760 3200 7812
rect 4344 7760 4396 7812
rect 4988 7760 5040 7812
rect 5356 7760 5408 7812
rect 5632 7828 5684 7880
rect 7472 7828 7524 7880
rect 9496 7828 9548 7880
rect 10692 7905 10701 7939
rect 10701 7905 10735 7939
rect 10735 7905 10744 7939
rect 10692 7896 10744 7905
rect 10784 7828 10836 7880
rect 12164 7871 12216 7880
rect 12164 7837 12173 7871
rect 12173 7837 12207 7871
rect 12207 7837 12216 7871
rect 12164 7828 12216 7837
rect 21364 8032 21416 8084
rect 9956 7760 10008 7812
rect 12716 7760 12768 7812
rect 13636 7803 13688 7812
rect 13636 7769 13654 7803
rect 13654 7769 13688 7803
rect 13636 7760 13688 7769
rect 15936 7871 15988 7880
rect 15936 7837 15945 7871
rect 15945 7837 15979 7871
rect 15979 7837 15988 7871
rect 15936 7828 15988 7837
rect 16028 7871 16080 7880
rect 16028 7837 16037 7871
rect 16037 7837 16071 7871
rect 16071 7837 16080 7871
rect 16028 7828 16080 7837
rect 16304 7803 16356 7812
rect 16304 7769 16338 7803
rect 16338 7769 16356 7803
rect 16304 7760 16356 7769
rect 7840 7692 7892 7744
rect 10324 7692 10376 7744
rect 12072 7735 12124 7744
rect 12072 7701 12081 7735
rect 12081 7701 12115 7735
rect 12115 7701 12124 7735
rect 12072 7692 12124 7701
rect 14188 7692 14240 7744
rect 14464 7692 14516 7744
rect 16120 7692 16172 7744
rect 17684 7760 17736 7812
rect 18512 7760 18564 7812
rect 18880 7871 18932 7880
rect 18880 7837 18889 7871
rect 18889 7837 18923 7871
rect 18923 7837 18932 7871
rect 18880 7828 18932 7837
rect 21824 7896 21876 7948
rect 18696 7692 18748 7744
rect 21548 7871 21600 7880
rect 21548 7837 21557 7871
rect 21557 7837 21591 7871
rect 21591 7837 21600 7871
rect 21548 7828 21600 7837
rect 21640 7828 21692 7880
rect 23020 7871 23072 7880
rect 23020 7837 23029 7871
rect 23029 7837 23063 7871
rect 23063 7837 23072 7871
rect 23020 7828 23072 7837
rect 23296 7871 23348 7880
rect 23296 7837 23305 7871
rect 23305 7837 23339 7871
rect 23339 7837 23348 7871
rect 23296 7828 23348 7837
rect 21732 7760 21784 7812
rect 22744 7803 22796 7812
rect 22744 7769 22762 7803
rect 22762 7769 22796 7803
rect 22744 7760 22796 7769
rect 21180 7692 21232 7744
rect 2658 7590 2710 7642
rect 2722 7590 2774 7642
rect 2786 7590 2838 7642
rect 2850 7590 2902 7642
rect 2914 7590 2966 7642
rect 2978 7590 3030 7642
rect 8658 7590 8710 7642
rect 8722 7590 8774 7642
rect 8786 7590 8838 7642
rect 8850 7590 8902 7642
rect 8914 7590 8966 7642
rect 8978 7590 9030 7642
rect 14658 7590 14710 7642
rect 14722 7590 14774 7642
rect 14786 7590 14838 7642
rect 14850 7590 14902 7642
rect 14914 7590 14966 7642
rect 14978 7590 15030 7642
rect 20658 7590 20710 7642
rect 20722 7590 20774 7642
rect 20786 7590 20838 7642
rect 20850 7590 20902 7642
rect 20914 7590 20966 7642
rect 20978 7590 21030 7642
rect 1676 7488 1728 7540
rect 2228 7488 2280 7540
rect 3792 7488 3844 7540
rect 3056 7420 3108 7472
rect 3148 7420 3200 7472
rect 3608 7463 3660 7472
rect 3608 7429 3620 7463
rect 3620 7429 3660 7463
rect 3608 7420 3660 7429
rect 4160 7420 4212 7472
rect 6092 7488 6144 7540
rect 7380 7488 7432 7540
rect 7840 7488 7892 7540
rect 6552 7420 6604 7472
rect 1952 7395 2004 7404
rect 1952 7361 1961 7395
rect 1961 7361 1995 7395
rect 1995 7361 2004 7395
rect 1952 7352 2004 7361
rect 4896 7352 4948 7404
rect 4988 7352 5040 7404
rect 5908 7395 5960 7404
rect 5908 7361 5926 7395
rect 5926 7361 5960 7395
rect 5908 7352 5960 7361
rect 6276 7352 6328 7404
rect 8392 7420 8444 7472
rect 9864 7531 9916 7540
rect 9864 7497 9873 7531
rect 9873 7497 9907 7531
rect 9907 7497 9916 7531
rect 9864 7488 9916 7497
rect 8208 7352 8260 7404
rect 8300 7352 8352 7404
rect 11336 7488 11388 7540
rect 11520 7420 11572 7472
rect 11796 7488 11848 7540
rect 13544 7531 13596 7540
rect 13544 7497 13553 7531
rect 13553 7497 13587 7531
rect 13587 7497 13596 7531
rect 13544 7488 13596 7497
rect 14280 7488 14332 7540
rect 15568 7488 15620 7540
rect 16764 7488 16816 7540
rect 21088 7488 21140 7540
rect 21272 7488 21324 7540
rect 21456 7531 21508 7540
rect 21456 7497 21465 7531
rect 21465 7497 21499 7531
rect 21499 7497 21508 7531
rect 21456 7488 21508 7497
rect 3056 7284 3108 7336
rect 3148 7284 3200 7336
rect 4436 7216 4488 7268
rect 6828 7284 6880 7336
rect 8392 7284 8444 7336
rect 11520 7284 11572 7336
rect 12072 7352 12124 7404
rect 12716 7352 12768 7404
rect 14372 7395 14424 7404
rect 14372 7361 14381 7395
rect 14381 7361 14415 7395
rect 14415 7361 14424 7395
rect 14372 7352 14424 7361
rect 15844 7395 15896 7404
rect 15844 7361 15862 7395
rect 15862 7361 15896 7395
rect 15844 7352 15896 7361
rect 11796 7284 11848 7336
rect 4620 7148 4672 7200
rect 5540 7148 5592 7200
rect 8116 7148 8168 7200
rect 8208 7148 8260 7200
rect 8392 7191 8444 7200
rect 8392 7157 8401 7191
rect 8401 7157 8435 7191
rect 8435 7157 8444 7191
rect 8392 7148 8444 7157
rect 11888 7259 11940 7268
rect 11888 7225 11897 7259
rect 11897 7225 11931 7259
rect 11931 7225 11940 7259
rect 11888 7216 11940 7225
rect 9864 7148 9916 7200
rect 9956 7191 10008 7200
rect 9956 7157 9965 7191
rect 9965 7157 9999 7191
rect 9999 7157 10008 7191
rect 9956 7148 10008 7157
rect 13452 7284 13504 7336
rect 13084 7148 13136 7200
rect 13544 7148 13596 7200
rect 18052 7327 18104 7336
rect 18052 7293 18061 7327
rect 18061 7293 18095 7327
rect 18095 7293 18104 7327
rect 18052 7284 18104 7293
rect 18328 7352 18380 7404
rect 19432 7352 19484 7404
rect 19708 7352 19760 7404
rect 19616 7327 19668 7336
rect 19616 7293 19625 7327
rect 19625 7293 19659 7327
rect 19659 7293 19668 7327
rect 19616 7284 19668 7293
rect 23296 7420 23348 7472
rect 21916 7352 21968 7404
rect 23112 7352 23164 7404
rect 21456 7216 21508 7268
rect 16948 7148 17000 7200
rect 23480 7148 23532 7200
rect 1918 7046 1970 7098
rect 1982 7046 2034 7098
rect 2046 7046 2098 7098
rect 2110 7046 2162 7098
rect 2174 7046 2226 7098
rect 2238 7046 2290 7098
rect 7918 7046 7970 7098
rect 7982 7046 8034 7098
rect 8046 7046 8098 7098
rect 8110 7046 8162 7098
rect 8174 7046 8226 7098
rect 8238 7046 8290 7098
rect 13918 7046 13970 7098
rect 13982 7046 14034 7098
rect 14046 7046 14098 7098
rect 14110 7046 14162 7098
rect 14174 7046 14226 7098
rect 14238 7046 14290 7098
rect 19918 7046 19970 7098
rect 19982 7046 20034 7098
rect 20046 7046 20098 7098
rect 20110 7046 20162 7098
rect 20174 7046 20226 7098
rect 20238 7046 20290 7098
rect 1308 6944 1360 6996
rect 1676 6944 1728 6996
rect 1768 6944 1820 6996
rect 2412 6944 2464 6996
rect 4160 6944 4212 6996
rect 1492 6808 1544 6860
rect 3056 6876 3108 6928
rect 4620 6944 4672 6996
rect 8392 6944 8444 6996
rect 10508 6944 10560 6996
rect 16304 6944 16356 6996
rect 18880 6944 18932 6996
rect 2780 6851 2832 6860
rect 2780 6817 2789 6851
rect 2789 6817 2823 6851
rect 2823 6817 2832 6851
rect 2780 6808 2832 6817
rect 2504 6740 2556 6792
rect 2872 6783 2924 6792
rect 2872 6749 2881 6783
rect 2881 6749 2915 6783
rect 2915 6749 2924 6783
rect 2872 6740 2924 6749
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 8300 6876 8352 6928
rect 9404 6876 9456 6928
rect 4252 6808 4304 6860
rect 8484 6808 8536 6860
rect 9496 6808 9548 6860
rect 19432 6944 19484 6996
rect 22008 6944 22060 6996
rect 22284 6944 22336 6996
rect 5816 6740 5868 6792
rect 7288 6783 7340 6792
rect 7288 6749 7297 6783
rect 7297 6749 7331 6783
rect 7331 6749 7340 6783
rect 7288 6740 7340 6749
rect 12440 6740 12492 6792
rect 13820 6740 13872 6792
rect 14096 6783 14148 6792
rect 14096 6749 14105 6783
rect 14105 6749 14139 6783
rect 14139 6749 14148 6783
rect 14096 6740 14148 6749
rect 14372 6783 14424 6792
rect 14372 6749 14406 6783
rect 14406 6749 14424 6783
rect 14372 6740 14424 6749
rect 18972 6740 19024 6792
rect 19248 6783 19300 6792
rect 19248 6749 19257 6783
rect 19257 6749 19291 6783
rect 19291 6749 19300 6783
rect 19248 6740 19300 6749
rect 21364 6740 21416 6792
rect 2688 6604 2740 6656
rect 7656 6672 7708 6724
rect 6276 6604 6328 6656
rect 6828 6604 6880 6656
rect 9680 6672 9732 6724
rect 9956 6672 10008 6724
rect 8484 6604 8536 6656
rect 11060 6604 11112 6656
rect 11244 6604 11296 6656
rect 13360 6604 13412 6656
rect 15752 6604 15804 6656
rect 17868 6672 17920 6724
rect 19524 6715 19576 6724
rect 19524 6681 19558 6715
rect 19558 6681 19576 6715
rect 19524 6672 19576 6681
rect 19708 6672 19760 6724
rect 22192 6808 22244 6860
rect 22928 6808 22980 6860
rect 17684 6604 17736 6656
rect 22560 6604 22612 6656
rect 2658 6502 2710 6554
rect 2722 6502 2774 6554
rect 2786 6502 2838 6554
rect 2850 6502 2902 6554
rect 2914 6502 2966 6554
rect 2978 6502 3030 6554
rect 8658 6502 8710 6554
rect 8722 6502 8774 6554
rect 8786 6502 8838 6554
rect 8850 6502 8902 6554
rect 8914 6502 8966 6554
rect 8978 6502 9030 6554
rect 14658 6502 14710 6554
rect 14722 6502 14774 6554
rect 14786 6502 14838 6554
rect 14850 6502 14902 6554
rect 14914 6502 14966 6554
rect 14978 6502 15030 6554
rect 20658 6502 20710 6554
rect 20722 6502 20774 6554
rect 20786 6502 20838 6554
rect 20850 6502 20902 6554
rect 20914 6502 20966 6554
rect 20978 6502 21030 6554
rect 1400 6400 1452 6452
rect 1584 6332 1636 6384
rect 4528 6332 4580 6384
rect 3056 6196 3108 6248
rect 4344 6264 4396 6316
rect 4620 6264 4672 6316
rect 4712 6264 4764 6316
rect 6184 6400 6236 6452
rect 6644 6400 6696 6452
rect 6920 6400 6972 6452
rect 7012 6400 7064 6452
rect 9864 6443 9916 6452
rect 9864 6409 9873 6443
rect 9873 6409 9907 6443
rect 9907 6409 9916 6443
rect 9864 6400 9916 6409
rect 10324 6400 10376 6452
rect 11336 6400 11388 6452
rect 7104 6264 7156 6316
rect 7564 6264 7616 6316
rect 9036 6264 9088 6316
rect 9496 6264 9548 6316
rect 9956 6307 10008 6316
rect 9956 6273 9965 6307
rect 9965 6273 9999 6307
rect 9999 6273 10008 6307
rect 9956 6264 10008 6273
rect 10232 6307 10284 6316
rect 10232 6273 10266 6307
rect 10266 6273 10284 6307
rect 10232 6264 10284 6273
rect 13636 6400 13688 6452
rect 15292 6400 15344 6452
rect 15936 6400 15988 6452
rect 16580 6400 16632 6452
rect 18512 6443 18564 6452
rect 18512 6409 18521 6443
rect 18521 6409 18555 6443
rect 18555 6409 18564 6443
rect 18512 6400 18564 6409
rect 18788 6400 18840 6452
rect 19248 6400 19300 6452
rect 23020 6400 23072 6452
rect 16672 6332 16724 6384
rect 13636 6307 13688 6316
rect 13636 6273 13654 6307
rect 13654 6273 13688 6307
rect 13636 6264 13688 6273
rect 13820 6264 13872 6316
rect 16120 6307 16172 6316
rect 16120 6273 16129 6307
rect 16129 6273 16163 6307
rect 16163 6273 16172 6307
rect 16120 6264 16172 6273
rect 16764 6264 16816 6316
rect 18144 6307 18196 6316
rect 18144 6273 18162 6307
rect 18162 6273 18196 6307
rect 18144 6264 18196 6273
rect 20996 6332 21048 6384
rect 19800 6264 19852 6316
rect 21180 6264 21232 6316
rect 21272 6264 21324 6316
rect 23112 6264 23164 6316
rect 23388 6264 23440 6316
rect 4344 6128 4396 6180
rect 6552 6196 6604 6248
rect 11704 6196 11756 6248
rect 14096 6239 14148 6248
rect 14096 6205 14105 6239
rect 14105 6205 14139 6239
rect 14139 6205 14148 6239
rect 14096 6196 14148 6205
rect 18420 6239 18472 6248
rect 18420 6205 18429 6239
rect 18429 6205 18463 6239
rect 18463 6205 18472 6239
rect 18420 6196 18472 6205
rect 4436 6060 4488 6112
rect 6644 6060 6696 6112
rect 11336 6103 11388 6112
rect 11336 6069 11345 6103
rect 11345 6069 11379 6103
rect 11379 6069 11388 6103
rect 11336 6060 11388 6069
rect 23204 6239 23256 6248
rect 23204 6205 23213 6239
rect 23213 6205 23247 6239
rect 23247 6205 23256 6239
rect 23204 6196 23256 6205
rect 14372 6060 14424 6112
rect 15476 6103 15528 6112
rect 15476 6069 15485 6103
rect 15485 6069 15519 6103
rect 15519 6069 15528 6103
rect 15476 6060 15528 6069
rect 15660 6060 15712 6112
rect 17040 6103 17092 6112
rect 17040 6069 17049 6103
rect 17049 6069 17083 6103
rect 17083 6069 17092 6103
rect 17040 6060 17092 6069
rect 20352 6060 20404 6112
rect 20904 6060 20956 6112
rect 1918 5958 1970 6010
rect 1982 5958 2034 6010
rect 2046 5958 2098 6010
rect 2110 5958 2162 6010
rect 2174 5958 2226 6010
rect 2238 5958 2290 6010
rect 7918 5958 7970 6010
rect 7982 5958 8034 6010
rect 8046 5958 8098 6010
rect 8110 5958 8162 6010
rect 8174 5958 8226 6010
rect 8238 5958 8290 6010
rect 13918 5958 13970 6010
rect 13982 5958 14034 6010
rect 14046 5958 14098 6010
rect 14110 5958 14162 6010
rect 14174 5958 14226 6010
rect 14238 5958 14290 6010
rect 19918 5958 19970 6010
rect 19982 5958 20034 6010
rect 20046 5958 20098 6010
rect 20110 5958 20162 6010
rect 20174 5958 20226 6010
rect 20238 5958 20290 6010
rect 1584 5856 1636 5908
rect 2780 5856 2832 5908
rect 3332 5856 3384 5908
rect 4068 5856 4120 5908
rect 4252 5856 4304 5908
rect 2504 5788 2556 5840
rect 3240 5788 3292 5840
rect 3792 5788 3844 5840
rect 1216 5652 1268 5704
rect 1952 5720 2004 5772
rect 2136 5695 2188 5704
rect 2136 5661 2145 5695
rect 2145 5661 2179 5695
rect 2179 5661 2188 5695
rect 2136 5652 2188 5661
rect 3056 5652 3108 5704
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 9128 5856 9180 5908
rect 10324 5856 10376 5908
rect 12716 5856 12768 5908
rect 12992 5856 13044 5908
rect 12624 5788 12676 5840
rect 13728 5788 13780 5840
rect 15660 5856 15712 5908
rect 18052 5856 18104 5908
rect 19616 5856 19668 5908
rect 20352 5856 20404 5908
rect 20904 5856 20956 5908
rect 20996 5899 21048 5908
rect 20996 5865 21005 5899
rect 21005 5865 21039 5899
rect 21039 5865 21048 5899
rect 20996 5856 21048 5865
rect 21548 5856 21600 5908
rect 22008 5899 22060 5908
rect 22008 5865 22017 5899
rect 22017 5865 22051 5899
rect 22051 5865 22060 5899
rect 22008 5856 22060 5865
rect 18144 5831 18196 5840
rect 18144 5797 18153 5831
rect 18153 5797 18187 5831
rect 18187 5797 18196 5831
rect 18144 5788 18196 5797
rect 19524 5831 19576 5840
rect 19524 5797 19533 5831
rect 19533 5797 19567 5831
rect 19567 5797 19576 5831
rect 19524 5788 19576 5797
rect 7196 5695 7248 5704
rect 7196 5661 7205 5695
rect 7205 5661 7239 5695
rect 7239 5661 7248 5695
rect 7196 5652 7248 5661
rect 8392 5652 8444 5704
rect 8484 5652 8536 5704
rect 3148 5584 3200 5636
rect 3516 5627 3568 5636
rect 3516 5593 3525 5627
rect 3525 5593 3559 5627
rect 3559 5593 3568 5627
rect 3516 5584 3568 5593
rect 4620 5627 4672 5636
rect 4620 5593 4632 5627
rect 4632 5593 4672 5627
rect 4620 5584 4672 5593
rect 4712 5584 4764 5636
rect 2412 5516 2464 5568
rect 3884 5516 3936 5568
rect 3976 5516 4028 5568
rect 5080 5516 5132 5568
rect 6460 5584 6512 5636
rect 6828 5516 6880 5568
rect 7380 5516 7432 5568
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 9220 5652 9272 5661
rect 9312 5695 9364 5704
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 17684 5720 17736 5772
rect 19340 5720 19392 5772
rect 9220 5516 9272 5568
rect 9496 5516 9548 5568
rect 10784 5695 10836 5704
rect 10784 5661 10793 5695
rect 10793 5661 10827 5695
rect 10827 5661 10836 5695
rect 10784 5652 10836 5661
rect 11060 5695 11112 5704
rect 11060 5661 11094 5695
rect 11094 5661 11112 5695
rect 11060 5652 11112 5661
rect 11336 5652 11388 5704
rect 10416 5584 10468 5636
rect 14188 5652 14240 5704
rect 11704 5516 11756 5568
rect 15660 5652 15712 5704
rect 16672 5695 16724 5704
rect 16672 5661 16681 5695
rect 16681 5661 16715 5695
rect 16715 5661 16724 5695
rect 16672 5652 16724 5661
rect 15108 5584 15160 5636
rect 15476 5584 15528 5636
rect 15384 5516 15436 5568
rect 18328 5652 18380 5704
rect 17408 5584 17460 5636
rect 19156 5652 19208 5704
rect 20168 5695 20220 5704
rect 20168 5661 20177 5695
rect 20177 5661 20211 5695
rect 20211 5661 20220 5695
rect 20168 5652 20220 5661
rect 21456 5720 21508 5772
rect 21824 5720 21876 5772
rect 21272 5584 21324 5636
rect 21640 5584 21692 5636
rect 23296 5695 23348 5704
rect 23296 5661 23305 5695
rect 23305 5661 23339 5695
rect 23339 5661 23348 5695
rect 23296 5652 23348 5661
rect 23388 5652 23440 5704
rect 18052 5559 18104 5568
rect 18052 5525 18061 5559
rect 18061 5525 18095 5559
rect 18095 5525 18104 5559
rect 18052 5516 18104 5525
rect 2658 5414 2710 5466
rect 2722 5414 2774 5466
rect 2786 5414 2838 5466
rect 2850 5414 2902 5466
rect 2914 5414 2966 5466
rect 2978 5414 3030 5466
rect 8658 5414 8710 5466
rect 8722 5414 8774 5466
rect 8786 5414 8838 5466
rect 8850 5414 8902 5466
rect 8914 5414 8966 5466
rect 8978 5414 9030 5466
rect 14658 5414 14710 5466
rect 14722 5414 14774 5466
rect 14786 5414 14838 5466
rect 14850 5414 14902 5466
rect 14914 5414 14966 5466
rect 14978 5414 15030 5466
rect 20658 5414 20710 5466
rect 20722 5414 20774 5466
rect 20786 5414 20838 5466
rect 20850 5414 20902 5466
rect 20914 5414 20966 5466
rect 20978 5414 21030 5466
rect 1952 5312 2004 5364
rect 2320 5312 2372 5364
rect 3700 5312 3752 5364
rect 3792 5312 3844 5364
rect 4620 5312 4672 5364
rect 7288 5312 7340 5364
rect 9036 5312 9088 5364
rect 9680 5312 9732 5364
rect 10048 5312 10100 5364
rect 13544 5312 13596 5364
rect 13820 5312 13872 5364
rect 14188 5312 14240 5364
rect 15292 5312 15344 5364
rect 15660 5355 15712 5364
rect 15660 5321 15669 5355
rect 15669 5321 15703 5355
rect 15703 5321 15712 5355
rect 15660 5312 15712 5321
rect 16028 5312 16080 5364
rect 17408 5355 17460 5364
rect 17408 5321 17417 5355
rect 17417 5321 17451 5355
rect 17451 5321 17460 5355
rect 17408 5312 17460 5321
rect 18420 5312 18472 5364
rect 19156 5312 19208 5364
rect 21272 5312 21324 5364
rect 21364 5355 21416 5364
rect 21364 5321 21373 5355
rect 21373 5321 21407 5355
rect 21407 5321 21416 5355
rect 21364 5312 21416 5321
rect 22376 5312 22428 5364
rect 23204 5312 23256 5364
rect 3976 5176 4028 5228
rect 4436 5176 4488 5228
rect 4896 5176 4948 5228
rect 6000 5219 6052 5228
rect 6000 5185 6009 5219
rect 6009 5185 6043 5219
rect 6043 5185 6052 5219
rect 6000 5176 6052 5185
rect 6460 5244 6512 5296
rect 10416 5244 10468 5296
rect 10508 5244 10560 5296
rect 12624 5244 12676 5296
rect 9404 5176 9456 5228
rect 9772 5176 9824 5228
rect 12900 5176 12952 5228
rect 14556 5176 14608 5228
rect 3516 5108 3568 5160
rect 7380 5108 7432 5160
rect 11336 5151 11388 5160
rect 11336 5117 11345 5151
rect 11345 5117 11379 5151
rect 11379 5117 11388 5151
rect 11336 5108 11388 5117
rect 13728 5151 13780 5160
rect 13728 5117 13737 5151
rect 13737 5117 13771 5151
rect 13771 5117 13780 5151
rect 13728 5108 13780 5117
rect 14464 5108 14516 5160
rect 15200 5176 15252 5228
rect 16948 5176 17000 5228
rect 18236 5176 18288 5228
rect 18328 5176 18380 5228
rect 19064 5176 19116 5228
rect 22468 5176 22520 5228
rect 23388 5176 23440 5228
rect 15844 5108 15896 5160
rect 19432 5108 19484 5160
rect 11704 5040 11756 5092
rect 7748 5015 7800 5024
rect 7748 4981 7757 5015
rect 7757 4981 7791 5015
rect 7791 4981 7800 5015
rect 7748 4972 7800 4981
rect 9680 5015 9732 5024
rect 9680 4981 9689 5015
rect 9689 4981 9723 5015
rect 9723 4981 9732 5015
rect 9680 4972 9732 4981
rect 10232 4972 10284 5024
rect 10692 4972 10744 5024
rect 12992 4972 13044 5024
rect 1918 4870 1970 4922
rect 1982 4870 2034 4922
rect 2046 4870 2098 4922
rect 2110 4870 2162 4922
rect 2174 4870 2226 4922
rect 2238 4870 2290 4922
rect 7918 4870 7970 4922
rect 7982 4870 8034 4922
rect 8046 4870 8098 4922
rect 8110 4870 8162 4922
rect 8174 4870 8226 4922
rect 8238 4870 8290 4922
rect 13918 4870 13970 4922
rect 13982 4870 14034 4922
rect 14046 4870 14098 4922
rect 14110 4870 14162 4922
rect 14174 4870 14226 4922
rect 14238 4870 14290 4922
rect 19918 4870 19970 4922
rect 19982 4870 20034 4922
rect 20046 4870 20098 4922
rect 20110 4870 20162 4922
rect 20174 4870 20226 4922
rect 20238 4870 20290 4922
rect 5816 4811 5868 4820
rect 5816 4777 5825 4811
rect 5825 4777 5859 4811
rect 5859 4777 5868 4811
rect 5816 4768 5868 4777
rect 7380 4768 7432 4820
rect 7564 4768 7616 4820
rect 9588 4768 9640 4820
rect 13084 4811 13136 4820
rect 13084 4777 13093 4811
rect 13093 4777 13127 4811
rect 13127 4777 13136 4811
rect 13084 4768 13136 4777
rect 13820 4768 13872 4820
rect 16672 4768 16724 4820
rect 17132 4768 17184 4820
rect 21732 4811 21784 4820
rect 21732 4777 21741 4811
rect 21741 4777 21775 4811
rect 21775 4777 21784 4811
rect 21732 4768 21784 4777
rect 22744 4768 22796 4820
rect 9404 4743 9456 4752
rect 9404 4709 9413 4743
rect 9413 4709 9447 4743
rect 9447 4709 9456 4743
rect 9404 4700 9456 4709
rect 4068 4632 4120 4684
rect 6000 4607 6052 4616
rect 6000 4573 6009 4607
rect 6009 4573 6043 4607
rect 6043 4573 6052 4607
rect 6000 4564 6052 4573
rect 6644 4607 6696 4616
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 6736 4564 6788 4616
rect 7104 4564 7156 4616
rect 7656 4564 7708 4616
rect 7748 4564 7800 4616
rect 8300 4564 8352 4616
rect 9036 4607 9088 4616
rect 9036 4573 9045 4607
rect 9045 4573 9079 4607
rect 9079 4573 9088 4607
rect 9036 4564 9088 4573
rect 9864 4632 9916 4684
rect 9956 4632 10008 4684
rect 8484 4496 8536 4548
rect 8116 4471 8168 4480
rect 8116 4437 8125 4471
rect 8125 4437 8159 4471
rect 8159 4437 8168 4471
rect 8116 4428 8168 4437
rect 11428 4607 11480 4616
rect 11428 4573 11437 4607
rect 11437 4573 11471 4607
rect 11471 4573 11480 4607
rect 11428 4564 11480 4573
rect 12992 4564 13044 4616
rect 13176 4607 13228 4616
rect 13176 4573 13185 4607
rect 13185 4573 13219 4607
rect 13219 4573 13228 4607
rect 13176 4564 13228 4573
rect 10048 4496 10100 4548
rect 10324 4496 10376 4548
rect 13544 4564 13596 4616
rect 22100 4632 22152 4684
rect 23480 4675 23532 4684
rect 23480 4641 23489 4675
rect 23489 4641 23523 4675
rect 23523 4641 23532 4675
rect 23480 4632 23532 4641
rect 14556 4564 14608 4616
rect 19064 4564 19116 4616
rect 9496 4428 9548 4480
rect 9588 4471 9640 4480
rect 9588 4437 9597 4471
rect 9597 4437 9631 4471
rect 9631 4437 9640 4471
rect 9588 4428 9640 4437
rect 12256 4428 12308 4480
rect 2658 4326 2710 4378
rect 2722 4326 2774 4378
rect 2786 4326 2838 4378
rect 2850 4326 2902 4378
rect 2914 4326 2966 4378
rect 2978 4326 3030 4378
rect 8658 4326 8710 4378
rect 8722 4326 8774 4378
rect 8786 4326 8838 4378
rect 8850 4326 8902 4378
rect 8914 4326 8966 4378
rect 8978 4326 9030 4378
rect 14658 4326 14710 4378
rect 14722 4326 14774 4378
rect 14786 4326 14838 4378
rect 14850 4326 14902 4378
rect 14914 4326 14966 4378
rect 14978 4326 15030 4378
rect 20658 4326 20710 4378
rect 20722 4326 20774 4378
rect 20786 4326 20838 4378
rect 20850 4326 20902 4378
rect 20914 4326 20966 4378
rect 20978 4326 21030 4378
rect 6000 4224 6052 4276
rect 8116 4224 8168 4276
rect 8300 4224 8352 4276
rect 9036 4224 9088 4276
rect 9772 4224 9824 4276
rect 13728 4224 13780 4276
rect 3424 4088 3476 4140
rect 6460 4131 6512 4140
rect 6460 4097 6469 4131
rect 6469 4097 6503 4131
rect 6503 4097 6512 4131
rect 6460 4088 6512 4097
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 6920 4088 6972 4140
rect 12624 4199 12676 4208
rect 12624 4165 12642 4199
rect 12642 4165 12676 4199
rect 12624 4156 12676 4165
rect 13176 4156 13228 4208
rect 8576 4088 8628 4140
rect 9864 4088 9916 4140
rect 9220 4020 9272 4072
rect 10784 4088 10836 4140
rect 11244 4088 11296 4140
rect 11888 4088 11940 4140
rect 10692 4063 10744 4072
rect 10692 4029 10701 4063
rect 10701 4029 10735 4063
rect 10735 4029 10744 4063
rect 10692 4020 10744 4029
rect 11060 3952 11112 4004
rect 22560 4131 22612 4140
rect 22560 4097 22569 4131
rect 22569 4097 22603 4131
rect 22603 4097 22612 4131
rect 22560 4088 22612 4097
rect 23112 4088 23164 4140
rect 14372 3952 14424 4004
rect 7288 3927 7340 3936
rect 7288 3893 7297 3927
rect 7297 3893 7331 3927
rect 7331 3893 7340 3927
rect 7288 3884 7340 3893
rect 8576 3884 8628 3936
rect 9128 3884 9180 3936
rect 12900 3884 12952 3936
rect 1918 3782 1970 3834
rect 1982 3782 2034 3834
rect 2046 3782 2098 3834
rect 2110 3782 2162 3834
rect 2174 3782 2226 3834
rect 2238 3782 2290 3834
rect 7918 3782 7970 3834
rect 7982 3782 8034 3834
rect 8046 3782 8098 3834
rect 8110 3782 8162 3834
rect 8174 3782 8226 3834
rect 8238 3782 8290 3834
rect 13918 3782 13970 3834
rect 13982 3782 14034 3834
rect 14046 3782 14098 3834
rect 14110 3782 14162 3834
rect 14174 3782 14226 3834
rect 14238 3782 14290 3834
rect 19918 3782 19970 3834
rect 19982 3782 20034 3834
rect 20046 3782 20098 3834
rect 20110 3782 20162 3834
rect 20174 3782 20226 3834
rect 20238 3782 20290 3834
rect 7196 3680 7248 3732
rect 8392 3680 8444 3732
rect 9036 3723 9088 3732
rect 9036 3689 9045 3723
rect 9045 3689 9079 3723
rect 9079 3689 9088 3723
rect 9036 3680 9088 3689
rect 9312 3680 9364 3732
rect 11336 3680 11388 3732
rect 12440 3723 12492 3732
rect 12440 3689 12449 3723
rect 12449 3689 12483 3723
rect 12483 3689 12492 3723
rect 12440 3680 12492 3689
rect 7472 3612 7524 3664
rect 8576 3612 8628 3664
rect 9404 3612 9456 3664
rect 11520 3655 11572 3664
rect 11520 3621 11529 3655
rect 11529 3621 11563 3655
rect 11563 3621 11572 3655
rect 11520 3612 11572 3621
rect 6460 3476 6512 3528
rect 8484 3476 8536 3528
rect 9496 3519 9548 3528
rect 9496 3485 9505 3519
rect 9505 3485 9539 3519
rect 9539 3485 9548 3519
rect 9496 3476 9548 3485
rect 9680 3476 9732 3528
rect 11060 3476 11112 3528
rect 11612 3476 11664 3528
rect 11980 3519 12032 3528
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 13544 3476 13596 3528
rect 2658 3238 2710 3290
rect 2722 3238 2774 3290
rect 2786 3238 2838 3290
rect 2850 3238 2902 3290
rect 2914 3238 2966 3290
rect 2978 3238 3030 3290
rect 8658 3238 8710 3290
rect 8722 3238 8774 3290
rect 8786 3238 8838 3290
rect 8850 3238 8902 3290
rect 8914 3238 8966 3290
rect 8978 3238 9030 3290
rect 14658 3238 14710 3290
rect 14722 3238 14774 3290
rect 14786 3238 14838 3290
rect 14850 3238 14902 3290
rect 14914 3238 14966 3290
rect 14978 3238 15030 3290
rect 20658 3238 20710 3290
rect 20722 3238 20774 3290
rect 20786 3238 20838 3290
rect 20850 3238 20902 3290
rect 20914 3238 20966 3290
rect 20978 3238 21030 3290
rect 6368 3000 6420 3052
rect 10968 2932 11020 2984
rect 1918 2694 1970 2746
rect 1982 2694 2034 2746
rect 2046 2694 2098 2746
rect 2110 2694 2162 2746
rect 2174 2694 2226 2746
rect 2238 2694 2290 2746
rect 7918 2694 7970 2746
rect 7982 2694 8034 2746
rect 8046 2694 8098 2746
rect 8110 2694 8162 2746
rect 8174 2694 8226 2746
rect 8238 2694 8290 2746
rect 13918 2694 13970 2746
rect 13982 2694 14034 2746
rect 14046 2694 14098 2746
rect 14110 2694 14162 2746
rect 14174 2694 14226 2746
rect 14238 2694 14290 2746
rect 19918 2694 19970 2746
rect 19982 2694 20034 2746
rect 20046 2694 20098 2746
rect 20110 2694 20162 2746
rect 20174 2694 20226 2746
rect 20238 2694 20290 2746
rect 6276 2524 6328 2576
rect 7196 2456 7248 2508
rect 5448 2388 5500 2440
rect 11796 2456 11848 2508
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 12256 2388 12308 2440
rect 12532 2431 12584 2440
rect 12532 2397 12541 2431
rect 12541 2397 12575 2431
rect 12575 2397 12584 2431
rect 12532 2388 12584 2397
rect 13360 2388 13412 2440
rect 17040 2388 17092 2440
rect 18236 2431 18288 2440
rect 18236 2397 18245 2431
rect 18245 2397 18279 2431
rect 18279 2397 18288 2431
rect 18236 2388 18288 2397
rect 7748 2320 7800 2372
rect 12164 2363 12216 2372
rect 12164 2329 12173 2363
rect 12173 2329 12207 2363
rect 12207 2329 12216 2363
rect 12164 2320 12216 2329
rect 12900 2320 12952 2372
rect 13544 2320 13596 2372
rect 17316 2363 17368 2372
rect 17316 2329 17325 2363
rect 17325 2329 17359 2363
rect 17359 2329 17368 2363
rect 17316 2320 17368 2329
rect 18052 2320 18104 2372
rect 2658 2150 2710 2202
rect 2722 2150 2774 2202
rect 2786 2150 2838 2202
rect 2850 2150 2902 2202
rect 2914 2150 2966 2202
rect 2978 2150 3030 2202
rect 8658 2150 8710 2202
rect 8722 2150 8774 2202
rect 8786 2150 8838 2202
rect 8850 2150 8902 2202
rect 8914 2150 8966 2202
rect 8978 2150 9030 2202
rect 14658 2150 14710 2202
rect 14722 2150 14774 2202
rect 14786 2150 14838 2202
rect 14850 2150 14902 2202
rect 14914 2150 14966 2202
rect 14978 2150 15030 2202
rect 20658 2150 20710 2202
rect 20722 2150 20774 2202
rect 20786 2150 20838 2202
rect 20850 2150 20902 2202
rect 20914 2150 20966 2202
rect 20978 2150 21030 2202
<< metal2 >>
rect 7746 26344 7802 27144
rect 8390 26344 8446 27144
rect 10966 26344 11022 27144
rect 13542 26344 13598 27144
rect 14186 26466 14242 27144
rect 14186 26438 14504 26466
rect 14186 26344 14242 26438
rect 1916 24508 2292 24517
rect 1972 24506 1996 24508
rect 2052 24506 2076 24508
rect 2132 24506 2156 24508
rect 2212 24506 2236 24508
rect 1972 24454 1982 24506
rect 2226 24454 2236 24506
rect 1972 24452 1996 24454
rect 2052 24452 2076 24454
rect 2132 24452 2156 24454
rect 2212 24452 2236 24454
rect 1916 24443 2292 24452
rect 7760 24274 7788 26344
rect 7916 24508 8292 24517
rect 7972 24506 7996 24508
rect 8052 24506 8076 24508
rect 8132 24506 8156 24508
rect 8212 24506 8236 24508
rect 7972 24454 7982 24506
rect 8226 24454 8236 24506
rect 7972 24452 7996 24454
rect 8052 24452 8076 24454
rect 8132 24452 8156 24454
rect 8212 24452 8236 24454
rect 7916 24443 8292 24452
rect 8404 24274 8432 26344
rect 10980 24274 11008 26344
rect 13556 24274 13584 26344
rect 13916 24508 14292 24517
rect 13972 24506 13996 24508
rect 14052 24506 14076 24508
rect 14132 24506 14156 24508
rect 14212 24506 14236 24508
rect 13972 24454 13982 24506
rect 14226 24454 14236 24506
rect 13972 24452 13996 24454
rect 14052 24452 14076 24454
rect 14132 24452 14156 24454
rect 14212 24452 14236 24454
rect 13916 24443 14292 24452
rect 14476 24274 14504 26438
rect 14830 26344 14886 27144
rect 14844 24274 14872 26344
rect 19916 24508 20292 24517
rect 19972 24506 19996 24508
rect 20052 24506 20076 24508
rect 20132 24506 20156 24508
rect 20212 24506 20236 24508
rect 19972 24454 19982 24506
rect 20226 24454 20236 24506
rect 19972 24452 19996 24454
rect 20052 24452 20076 24454
rect 20132 24452 20156 24454
rect 20212 24452 20236 24454
rect 19916 24443 20292 24452
rect 7748 24268 7800 24274
rect 7748 24210 7800 24216
rect 8392 24268 8444 24274
rect 8392 24210 8444 24216
rect 10968 24268 11020 24274
rect 10968 24210 11020 24216
rect 13544 24268 13596 24274
rect 13544 24210 13596 24216
rect 14464 24268 14516 24274
rect 14464 24210 14516 24216
rect 14832 24268 14884 24274
rect 14832 24210 14884 24216
rect 7564 24200 7616 24206
rect 7564 24142 7616 24148
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 10784 24200 10836 24206
rect 10784 24142 10836 24148
rect 12992 24200 13044 24206
rect 12992 24142 13044 24148
rect 14556 24200 14608 24206
rect 14556 24142 14608 24148
rect 15384 24200 15436 24206
rect 15384 24142 15436 24148
rect 2656 23964 3032 23973
rect 2712 23962 2736 23964
rect 2792 23962 2816 23964
rect 2872 23962 2896 23964
rect 2952 23962 2976 23964
rect 2712 23910 2722 23962
rect 2966 23910 2976 23962
rect 2712 23908 2736 23910
rect 2792 23908 2816 23910
rect 2872 23908 2896 23910
rect 2952 23908 2976 23910
rect 2656 23899 3032 23908
rect 1916 23420 2292 23429
rect 1972 23418 1996 23420
rect 2052 23418 2076 23420
rect 2132 23418 2156 23420
rect 2212 23418 2236 23420
rect 1972 23366 1982 23418
rect 2226 23366 2236 23418
rect 1972 23364 1996 23366
rect 2052 23364 2076 23366
rect 2132 23364 2156 23366
rect 2212 23364 2236 23366
rect 1916 23355 2292 23364
rect 2656 22876 3032 22885
rect 2712 22874 2736 22876
rect 2792 22874 2816 22876
rect 2872 22874 2896 22876
rect 2952 22874 2976 22876
rect 2712 22822 2722 22874
rect 2966 22822 2976 22874
rect 2712 22820 2736 22822
rect 2792 22820 2816 22822
rect 2872 22820 2896 22822
rect 2952 22820 2976 22822
rect 2656 22811 3032 22820
rect 1916 22332 2292 22341
rect 1972 22330 1996 22332
rect 2052 22330 2076 22332
rect 2132 22330 2156 22332
rect 2212 22330 2236 22332
rect 1972 22278 1982 22330
rect 2226 22278 2236 22330
rect 1972 22276 1996 22278
rect 2052 22276 2076 22278
rect 2132 22276 2156 22278
rect 2212 22276 2236 22278
rect 1916 22267 2292 22276
rect 6828 21888 6880 21894
rect 6828 21830 6880 21836
rect 2656 21788 3032 21797
rect 2712 21786 2736 21788
rect 2792 21786 2816 21788
rect 2872 21786 2896 21788
rect 2952 21786 2976 21788
rect 2712 21734 2722 21786
rect 2966 21734 2976 21786
rect 2712 21732 2736 21734
rect 2792 21732 2816 21734
rect 2872 21732 2896 21734
rect 2952 21732 2976 21734
rect 2656 21723 3032 21732
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 1916 21244 2292 21253
rect 1972 21242 1996 21244
rect 2052 21242 2076 21244
rect 2132 21242 2156 21244
rect 2212 21242 2236 21244
rect 1972 21190 1982 21242
rect 2226 21190 2236 21242
rect 1972 21188 1996 21190
rect 2052 21188 2076 21190
rect 2132 21188 2156 21190
rect 2212 21188 2236 21190
rect 1916 21179 2292 21188
rect 5540 21004 5592 21010
rect 5540 20946 5592 20952
rect 4896 20868 4948 20874
rect 4896 20810 4948 20816
rect 4344 20800 4396 20806
rect 4344 20742 4396 20748
rect 2656 20700 3032 20709
rect 2712 20698 2736 20700
rect 2792 20698 2816 20700
rect 2872 20698 2896 20700
rect 2952 20698 2976 20700
rect 2712 20646 2722 20698
rect 2966 20646 2976 20698
rect 2712 20644 2736 20646
rect 2792 20644 2816 20646
rect 2872 20644 2896 20646
rect 2952 20644 2976 20646
rect 2656 20635 3032 20644
rect 1916 20156 2292 20165
rect 1972 20154 1996 20156
rect 2052 20154 2076 20156
rect 2132 20154 2156 20156
rect 2212 20154 2236 20156
rect 1972 20102 1982 20154
rect 2226 20102 2236 20154
rect 1972 20100 1996 20102
rect 2052 20100 2076 20102
rect 2132 20100 2156 20102
rect 2212 20100 2236 20102
rect 1916 20091 2292 20100
rect 3790 19816 3846 19825
rect 3790 19751 3846 19760
rect 2656 19612 3032 19621
rect 2712 19610 2736 19612
rect 2792 19610 2816 19612
rect 2872 19610 2896 19612
rect 2952 19610 2976 19612
rect 2712 19558 2722 19610
rect 2966 19558 2976 19610
rect 2712 19556 2736 19558
rect 2792 19556 2816 19558
rect 2872 19556 2896 19558
rect 2952 19556 2976 19558
rect 2656 19547 3032 19556
rect 1916 19068 2292 19077
rect 1972 19066 1996 19068
rect 2052 19066 2076 19068
rect 2132 19066 2156 19068
rect 2212 19066 2236 19068
rect 1972 19014 1982 19066
rect 2226 19014 2236 19066
rect 1972 19012 1996 19014
rect 2052 19012 2076 19014
rect 2132 19012 2156 19014
rect 2212 19012 2236 19014
rect 1916 19003 2292 19012
rect 2656 18524 3032 18533
rect 2712 18522 2736 18524
rect 2792 18522 2816 18524
rect 2872 18522 2896 18524
rect 2952 18522 2976 18524
rect 2712 18470 2722 18522
rect 2966 18470 2976 18522
rect 2712 18468 2736 18470
rect 2792 18468 2816 18470
rect 2872 18468 2896 18470
rect 2952 18468 2976 18470
rect 2656 18459 3032 18468
rect 1916 17980 2292 17989
rect 1972 17978 1996 17980
rect 2052 17978 2076 17980
rect 2132 17978 2156 17980
rect 2212 17978 2236 17980
rect 1972 17926 1982 17978
rect 2226 17926 2236 17978
rect 1972 17924 1996 17926
rect 2052 17924 2076 17926
rect 2132 17924 2156 17926
rect 2212 17924 2236 17926
rect 1916 17915 2292 17924
rect 3516 17536 3568 17542
rect 3516 17478 3568 17484
rect 2656 17436 3032 17445
rect 2712 17434 2736 17436
rect 2792 17434 2816 17436
rect 2872 17434 2896 17436
rect 2952 17434 2976 17436
rect 2712 17382 2722 17434
rect 2966 17382 2976 17434
rect 2712 17380 2736 17382
rect 2792 17380 2816 17382
rect 2872 17380 2896 17382
rect 2952 17380 2976 17382
rect 2656 17371 3032 17380
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 940 17128 992 17134
rect 938 17096 940 17105
rect 992 17096 994 17105
rect 938 17031 994 17040
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 1916 16892 2292 16901
rect 1972 16890 1996 16892
rect 2052 16890 2076 16892
rect 2132 16890 2156 16892
rect 2212 16890 2236 16892
rect 1972 16838 1982 16890
rect 2226 16838 2236 16890
rect 1972 16836 1996 16838
rect 2052 16836 2076 16838
rect 2132 16836 2156 16838
rect 2212 16836 2236 16838
rect 1916 16827 2292 16836
rect 2136 16584 2188 16590
rect 2136 16526 2188 16532
rect 1216 16448 1268 16454
rect 1216 16390 1268 16396
rect 940 16040 992 16046
rect 940 15982 992 15988
rect 952 15745 980 15982
rect 938 15736 994 15745
rect 938 15671 994 15680
rect 938 13696 994 13705
rect 938 13631 994 13640
rect 952 13394 980 13631
rect 940 13388 992 13394
rect 940 13330 992 13336
rect 938 12336 994 12345
rect 938 12271 994 12280
rect 952 12238 980 12271
rect 940 12232 992 12238
rect 940 12174 992 12180
rect 1228 10674 1256 16390
rect 1492 16176 1544 16182
rect 1492 16118 1544 16124
rect 1308 14340 1360 14346
rect 1308 14282 1360 14288
rect 1320 13161 1348 14282
rect 1504 13682 1532 16118
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1676 16040 1728 16046
rect 1872 16017 1900 16050
rect 1676 15982 1728 15988
rect 1858 16008 1914 16017
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1596 15162 1624 15302
rect 1584 15156 1636 15162
rect 1584 15098 1636 15104
rect 1688 14906 1716 15982
rect 2148 15994 2176 16526
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2148 15966 2360 15994
rect 1858 15943 1914 15952
rect 1916 15804 2292 15813
rect 1972 15802 1996 15804
rect 2052 15802 2076 15804
rect 2132 15802 2156 15804
rect 2212 15802 2236 15804
rect 1972 15750 1982 15802
rect 2226 15750 2236 15802
rect 1972 15748 1996 15750
rect 2052 15748 2076 15750
rect 2132 15748 2156 15750
rect 2212 15748 2236 15750
rect 1916 15739 2292 15748
rect 2226 15600 2282 15609
rect 2226 15535 2282 15544
rect 2240 15502 2268 15535
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 1860 15428 1912 15434
rect 1860 15370 1912 15376
rect 1768 15360 1820 15366
rect 1768 15302 1820 15308
rect 1596 14878 1716 14906
rect 1596 14464 1624 14878
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1688 14618 1716 14758
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1596 14436 1716 14464
rect 1504 13654 1624 13682
rect 1306 13152 1362 13161
rect 1306 13087 1362 13096
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1216 10668 1268 10674
rect 1216 10610 1268 10616
rect 1308 9920 1360 9926
rect 1308 9862 1360 9868
rect 1214 7984 1270 7993
rect 1214 7919 1270 7928
rect 1228 5710 1256 7919
rect 1320 7002 1348 9862
rect 1308 6996 1360 7002
rect 1308 6938 1360 6944
rect 1412 6458 1440 12242
rect 1596 11898 1624 13654
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1504 6866 1532 11630
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1596 6390 1624 10202
rect 1688 7857 1716 14436
rect 1780 13938 1808 15302
rect 1872 14958 1900 15370
rect 2136 15360 2188 15366
rect 2136 15302 2188 15308
rect 1860 14952 1912 14958
rect 1860 14894 1912 14900
rect 2148 14822 2176 15302
rect 2136 14816 2188 14822
rect 2136 14758 2188 14764
rect 1916 14716 2292 14725
rect 1972 14714 1996 14716
rect 2052 14714 2076 14716
rect 2132 14714 2156 14716
rect 2212 14714 2236 14716
rect 1972 14662 1982 14714
rect 2226 14662 2236 14714
rect 1972 14660 1996 14662
rect 2052 14660 2076 14662
rect 2132 14660 2156 14662
rect 2212 14660 2236 14662
rect 1916 14651 2292 14660
rect 2136 14340 2188 14346
rect 2136 14282 2188 14288
rect 2148 13938 2176 14282
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 1916 13628 2292 13637
rect 1972 13626 1996 13628
rect 2052 13626 2076 13628
rect 2132 13626 2156 13628
rect 2212 13626 2236 13628
rect 1972 13574 1982 13626
rect 2226 13574 2236 13626
rect 1972 13572 1996 13574
rect 2052 13572 2076 13574
rect 2132 13572 2156 13574
rect 2212 13572 2236 13574
rect 1916 13563 2292 13572
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1780 11830 1808 12582
rect 1916 12540 2292 12549
rect 1972 12538 1996 12540
rect 2052 12538 2076 12540
rect 2132 12538 2156 12540
rect 2212 12538 2236 12540
rect 1972 12486 1982 12538
rect 2226 12486 2236 12538
rect 1972 12484 1996 12486
rect 2052 12484 2076 12486
rect 2132 12484 2156 12486
rect 2212 12484 2236 12486
rect 1916 12475 2292 12484
rect 1768 11824 1820 11830
rect 1768 11766 1820 11772
rect 1766 11656 1822 11665
rect 1766 11591 1768 11600
rect 1820 11591 1822 11600
rect 1768 11562 1820 11568
rect 1916 11452 2292 11461
rect 1972 11450 1996 11452
rect 2052 11450 2076 11452
rect 2132 11450 2156 11452
rect 2212 11450 2236 11452
rect 1972 11398 1982 11450
rect 2226 11398 2236 11450
rect 1972 11396 1996 11398
rect 2052 11396 2076 11398
rect 2132 11396 2156 11398
rect 2212 11396 2236 11398
rect 1916 11387 2292 11396
rect 2332 11234 2360 15966
rect 2424 15366 2452 16390
rect 2656 16348 3032 16357
rect 2712 16346 2736 16348
rect 2792 16346 2816 16348
rect 2872 16346 2896 16348
rect 2952 16346 2976 16348
rect 2712 16294 2722 16346
rect 2966 16294 2976 16346
rect 2712 16292 2736 16294
rect 2792 16292 2816 16294
rect 2872 16292 2896 16294
rect 2952 16292 2976 16294
rect 2656 16283 3032 16292
rect 2504 16040 2556 16046
rect 2556 15988 2636 15994
rect 2504 15982 2636 15988
rect 2516 15966 2636 15982
rect 2504 15904 2556 15910
rect 2504 15846 2556 15852
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2240 11206 2360 11234
rect 2240 10742 2268 11206
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2228 10736 2280 10742
rect 2228 10678 2280 10684
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1872 10554 1900 10610
rect 1780 10526 1900 10554
rect 1674 7848 1730 7857
rect 1674 7783 1730 7792
rect 1688 7546 1716 7783
rect 1780 7698 1808 10526
rect 1916 10364 2292 10373
rect 1972 10362 1996 10364
rect 2052 10362 2076 10364
rect 2132 10362 2156 10364
rect 2212 10362 2236 10364
rect 1972 10310 1982 10362
rect 2226 10310 2236 10362
rect 1972 10308 1996 10310
rect 2052 10308 2076 10310
rect 2132 10308 2156 10310
rect 2212 10308 2236 10310
rect 1916 10299 2292 10308
rect 2228 10056 2280 10062
rect 2228 9998 2280 10004
rect 2240 9722 2268 9998
rect 2228 9716 2280 9722
rect 2228 9658 2280 9664
rect 2226 9616 2282 9625
rect 2226 9551 2228 9560
rect 2280 9551 2282 9560
rect 2228 9522 2280 9528
rect 1916 9276 2292 9285
rect 1972 9274 1996 9276
rect 2052 9274 2076 9276
rect 2132 9274 2156 9276
rect 2212 9274 2236 9276
rect 1972 9222 1982 9274
rect 2226 9222 2236 9274
rect 1972 9220 1996 9222
rect 2052 9220 2076 9222
rect 2132 9220 2156 9222
rect 2212 9220 2236 9222
rect 1916 9211 2292 9220
rect 2332 9160 2360 11086
rect 2424 9674 2452 15302
rect 2516 11830 2544 15846
rect 2608 15473 2636 15966
rect 2594 15464 2650 15473
rect 2594 15399 2650 15408
rect 2656 15260 3032 15269
rect 2712 15258 2736 15260
rect 2792 15258 2816 15260
rect 2872 15258 2896 15260
rect 2952 15258 2976 15260
rect 2712 15206 2722 15258
rect 2966 15206 2976 15258
rect 2712 15204 2736 15206
rect 2792 15204 2816 15206
rect 2872 15204 2896 15206
rect 2952 15204 2976 15206
rect 2656 15195 3032 15204
rect 3068 15094 3096 16934
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3252 15162 3280 16594
rect 3344 16250 3372 17138
rect 3436 17105 3464 17138
rect 3422 17096 3478 17105
rect 3422 17031 3478 17040
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3436 16182 3464 16390
rect 3424 16176 3476 16182
rect 3424 16118 3476 16124
rect 3528 15570 3556 17478
rect 3700 16244 3752 16250
rect 3700 16186 3752 16192
rect 3606 16144 3662 16153
rect 3712 16114 3740 16186
rect 3606 16079 3662 16088
rect 3700 16108 3752 16114
rect 3620 16046 3648 16079
rect 3700 16050 3752 16056
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3606 15600 3662 15609
rect 3516 15564 3568 15570
rect 3606 15535 3662 15544
rect 3516 15506 3568 15512
rect 3620 15502 3648 15535
rect 3712 15502 3740 15846
rect 3608 15496 3660 15502
rect 3608 15438 3660 15444
rect 3700 15496 3752 15502
rect 3700 15438 3752 15444
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 3056 15088 3108 15094
rect 3056 15030 3108 15036
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2608 14346 2636 14758
rect 2596 14340 2648 14346
rect 2596 14282 2648 14288
rect 2656 14172 3032 14181
rect 2712 14170 2736 14172
rect 2792 14170 2816 14172
rect 2872 14170 2896 14172
rect 2952 14170 2976 14172
rect 2712 14118 2722 14170
rect 2966 14118 2976 14170
rect 2712 14116 2736 14118
rect 2792 14116 2816 14118
rect 2872 14116 2896 14118
rect 2952 14116 2976 14118
rect 2656 14107 3032 14116
rect 3160 13938 3188 14962
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 3068 13326 3096 13670
rect 3252 13530 3280 15098
rect 3344 14482 3372 15302
rect 3700 15088 3752 15094
rect 3700 15030 3752 15036
rect 3712 14906 3740 15030
rect 3528 14878 3740 14906
rect 3528 14550 3556 14878
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3620 14550 3648 14758
rect 3516 14544 3568 14550
rect 3516 14486 3568 14492
rect 3608 14544 3660 14550
rect 3608 14486 3660 14492
rect 3332 14476 3384 14482
rect 3332 14418 3384 14424
rect 3424 14340 3476 14346
rect 3424 14282 3476 14288
rect 3436 14226 3464 14282
rect 3700 14272 3752 14278
rect 3436 14220 3700 14226
rect 3436 14214 3752 14220
rect 3436 14198 3740 14214
rect 3700 14000 3752 14006
rect 3700 13942 3752 13948
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 3344 13410 3372 13874
rect 3344 13382 3556 13410
rect 3528 13326 3556 13382
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 3516 13320 3568 13326
rect 3712 13308 3740 13942
rect 3804 13433 3832 19751
rect 4356 19334 4384 20742
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 4816 19378 4844 20402
rect 4172 19306 4384 19334
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 3884 18760 3936 18766
rect 3884 18702 3936 18708
rect 3896 18426 3924 18702
rect 3884 18420 3936 18426
rect 3884 18362 3936 18368
rect 4172 18290 4200 19306
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 4540 18766 4568 19110
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 4632 18698 4660 19314
rect 4620 18692 4672 18698
rect 4620 18634 4672 18640
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 4172 17542 4200 18226
rect 4712 17808 4764 17814
rect 4712 17750 4764 17756
rect 4252 17740 4304 17746
rect 4252 17682 4304 17688
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 4264 17202 4292 17682
rect 4724 17338 4752 17750
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4528 17264 4580 17270
rect 4528 17206 4580 17212
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4436 17196 4488 17202
rect 4436 17138 4488 17144
rect 3882 16688 3938 16697
rect 3882 16623 3938 16632
rect 3896 15706 3924 16623
rect 3884 15700 3936 15706
rect 3884 15642 3936 15648
rect 3988 15502 4016 17138
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4160 16516 4212 16522
rect 4160 16458 4212 16464
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4080 16182 4108 16390
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 4068 15632 4120 15638
rect 4068 15574 4120 15580
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3884 14340 3936 14346
rect 3884 14282 3936 14288
rect 3896 13938 3924 14282
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3790 13424 3846 13433
rect 4080 13394 4108 15574
rect 4172 15026 4200 16458
rect 4264 15570 4292 16934
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4250 15464 4306 15473
rect 4250 15399 4306 15408
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 3790 13359 3846 13368
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 3712 13280 3832 13308
rect 3516 13262 3568 13268
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 3332 13252 3384 13258
rect 3332 13194 3384 13200
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 2656 13084 3032 13093
rect 2712 13082 2736 13084
rect 2792 13082 2816 13084
rect 2872 13082 2896 13084
rect 2952 13082 2976 13084
rect 2712 13030 2722 13082
rect 2966 13030 2976 13082
rect 2712 13028 2736 13030
rect 2792 13028 2816 13030
rect 2872 13028 2896 13030
rect 2952 13028 2976 13030
rect 2656 13019 3032 13028
rect 3160 12918 3188 13126
rect 3148 12912 3200 12918
rect 3148 12854 3200 12860
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2976 12434 3004 12786
rect 2976 12406 3188 12434
rect 2656 11996 3032 12005
rect 2712 11994 2736 11996
rect 2792 11994 2816 11996
rect 2872 11994 2896 11996
rect 2952 11994 2976 11996
rect 2712 11942 2722 11994
rect 2966 11942 2976 11994
rect 2712 11940 2736 11942
rect 2792 11940 2816 11942
rect 2872 11940 2896 11942
rect 2952 11940 2976 11942
rect 2656 11931 3032 11940
rect 2504 11824 2556 11830
rect 2504 11766 2556 11772
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 2656 10908 3032 10917
rect 2712 10906 2736 10908
rect 2792 10906 2816 10908
rect 2872 10906 2896 10908
rect 2952 10906 2976 10908
rect 2712 10854 2722 10906
rect 2966 10854 2976 10906
rect 2712 10852 2736 10854
rect 2792 10852 2816 10854
rect 2872 10852 2896 10854
rect 2952 10852 2976 10854
rect 2656 10843 3032 10852
rect 2504 10736 2556 10742
rect 2504 10678 2556 10684
rect 2516 10266 2544 10678
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2608 10062 2636 10610
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2656 9820 3032 9829
rect 2712 9818 2736 9820
rect 2792 9818 2816 9820
rect 2872 9818 2896 9820
rect 2952 9818 2976 9820
rect 2712 9766 2722 9818
rect 2966 9766 2976 9818
rect 2712 9764 2736 9766
rect 2792 9764 2816 9766
rect 2872 9764 2896 9766
rect 2952 9764 2976 9766
rect 2656 9755 3032 9764
rect 2424 9646 2636 9674
rect 2410 9480 2466 9489
rect 2608 9450 2636 9646
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2596 9444 2648 9450
rect 2410 9415 2412 9424
rect 2464 9415 2466 9424
rect 2412 9386 2464 9392
rect 2516 9404 2596 9432
rect 2056 9132 2360 9160
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1872 8498 1900 8842
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 2056 8276 2084 9132
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2148 8498 2176 8910
rect 2516 8650 2544 9404
rect 2596 9386 2648 9392
rect 2976 8974 3004 9454
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2656 8732 3032 8741
rect 2712 8730 2736 8732
rect 2792 8730 2816 8732
rect 2872 8730 2896 8732
rect 2952 8730 2976 8732
rect 2712 8678 2722 8730
rect 2966 8678 2976 8730
rect 2712 8676 2736 8678
rect 2792 8676 2816 8678
rect 2872 8676 2896 8678
rect 2952 8676 2976 8678
rect 2656 8667 3032 8676
rect 2424 8622 2544 8650
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2056 8248 2360 8276
rect 1916 8188 2292 8197
rect 1972 8186 1996 8188
rect 2052 8186 2076 8188
rect 2132 8186 2156 8188
rect 2212 8186 2236 8188
rect 1972 8134 1982 8186
rect 2226 8134 2236 8186
rect 1972 8132 1996 8134
rect 2052 8132 2076 8134
rect 2132 8132 2156 8134
rect 2212 8132 2236 8134
rect 1916 8123 2292 8132
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 1780 7670 1900 7698
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1872 7256 1900 7670
rect 2240 7546 2268 8026
rect 2332 7970 2360 8248
rect 2424 8090 2452 8622
rect 2504 8560 2556 8566
rect 2504 8502 2556 8508
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2332 7942 2452 7970
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1688 7228 1900 7256
rect 1688 7002 1716 7228
rect 1964 7188 1992 7346
rect 1780 7160 1992 7188
rect 1780 7002 1808 7160
rect 1916 7100 2292 7109
rect 1972 7098 1996 7100
rect 2052 7098 2076 7100
rect 2132 7098 2156 7100
rect 2212 7098 2236 7100
rect 1972 7046 1982 7098
rect 2226 7046 2236 7098
rect 1972 7044 1996 7046
rect 2052 7044 2076 7046
rect 2132 7044 2156 7046
rect 2212 7044 2236 7046
rect 1916 7035 2292 7044
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1584 6384 1636 6390
rect 1584 6326 1636 6332
rect 1596 5914 1624 6326
rect 1916 6012 2292 6021
rect 1972 6010 1996 6012
rect 2052 6010 2076 6012
rect 2132 6010 2156 6012
rect 2212 6010 2236 6012
rect 1972 5958 1982 6010
rect 2226 5958 2236 6010
rect 1972 5956 1996 5958
rect 2052 5956 2076 5958
rect 2132 5956 2156 5958
rect 2212 5956 2236 5958
rect 1916 5947 2292 5956
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 2226 5808 2282 5817
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 2148 5766 2226 5794
rect 1216 5704 1268 5710
rect 1216 5646 1268 5652
rect 1964 5370 1992 5714
rect 2148 5710 2176 5766
rect 2226 5743 2282 5752
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 2332 5370 2360 7822
rect 2424 7002 2452 7942
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2516 6798 2544 8502
rect 2594 7984 2650 7993
rect 2594 7919 2650 7928
rect 2608 7818 2636 7919
rect 2596 7812 2648 7818
rect 2596 7754 2648 7760
rect 2656 7644 3032 7653
rect 2712 7642 2736 7644
rect 2792 7642 2816 7644
rect 2872 7642 2896 7644
rect 2952 7642 2976 7644
rect 2712 7590 2722 7642
rect 2966 7590 2976 7642
rect 2712 7588 2736 7590
rect 2792 7588 2816 7590
rect 2872 7588 2896 7590
rect 2952 7588 2976 7590
rect 2656 7579 3032 7588
rect 3068 7478 3096 11630
rect 3160 10674 3188 12406
rect 3252 11762 3280 13194
rect 3344 12442 3372 13194
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3332 12436 3384 12442
rect 3436 12434 3464 12786
rect 3528 12646 3556 13262
rect 3804 12889 3832 13280
rect 3790 12880 3846 12889
rect 3790 12815 3846 12824
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3436 12406 3556 12434
rect 3332 12378 3384 12384
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3344 11558 3372 12174
rect 3528 11558 3556 12406
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3344 11218 3372 11494
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3252 9382 3280 11018
rect 3332 10668 3384 10674
rect 3384 10628 3464 10656
rect 3332 10610 3384 10616
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3344 8566 3372 9590
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3148 7812 3200 7818
rect 3148 7754 3200 7760
rect 3160 7478 3188 7754
rect 3056 7472 3108 7478
rect 3056 7414 3108 7420
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3056 7336 3108 7342
rect 3054 7304 3056 7313
rect 3148 7336 3200 7342
rect 3108 7304 3110 7313
rect 3148 7278 3200 7284
rect 3054 7239 3110 7248
rect 2686 7168 2742 7177
rect 2686 7103 2742 7112
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2410 6080 2466 6089
rect 2410 6015 2466 6024
rect 2424 5574 2452 6015
rect 2516 5846 2544 6734
rect 2700 6662 2728 7103
rect 2778 7032 2834 7041
rect 2778 6967 2834 6976
rect 2792 6866 2820 6967
rect 3056 6928 3108 6934
rect 3054 6896 3056 6905
rect 3108 6896 3110 6905
rect 2780 6860 2832 6866
rect 3054 6831 3110 6840
rect 2780 6802 2832 6808
rect 2872 6792 2924 6798
rect 2924 6752 3096 6780
rect 2872 6734 2924 6740
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2656 6556 3032 6565
rect 2712 6554 2736 6556
rect 2792 6554 2816 6556
rect 2872 6554 2896 6556
rect 2952 6554 2976 6556
rect 2712 6502 2722 6554
rect 2966 6502 2976 6554
rect 2712 6500 2736 6502
rect 2792 6500 2816 6502
rect 2872 6500 2896 6502
rect 2952 6500 2976 6502
rect 2656 6491 3032 6500
rect 3068 6361 3096 6752
rect 3054 6352 3110 6361
rect 3054 6287 3110 6296
rect 3056 6248 3108 6254
rect 3054 6216 3056 6225
rect 3108 6216 3110 6225
rect 3054 6151 3110 6160
rect 3054 5944 3110 5953
rect 2780 5908 2832 5914
rect 3054 5879 3110 5888
rect 2780 5850 2832 5856
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 2792 5658 2820 5850
rect 3068 5710 3096 5879
rect 3056 5704 3108 5710
rect 2870 5672 2926 5681
rect 2792 5630 2870 5658
rect 3056 5646 3108 5652
rect 3160 5642 3188 7278
rect 3252 5846 3280 8366
rect 3344 5914 3372 8366
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 2870 5607 2926 5616
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2656 5468 3032 5477
rect 2712 5466 2736 5468
rect 2792 5466 2816 5468
rect 2872 5466 2896 5468
rect 2952 5466 2976 5468
rect 2712 5414 2722 5466
rect 2966 5414 2976 5466
rect 2712 5412 2736 5414
rect 2792 5412 2816 5414
rect 2872 5412 2896 5414
rect 2952 5412 2976 5414
rect 2656 5403 3032 5412
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 1916 4924 2292 4933
rect 1972 4922 1996 4924
rect 2052 4922 2076 4924
rect 2132 4922 2156 4924
rect 2212 4922 2236 4924
rect 1972 4870 1982 4922
rect 2226 4870 2236 4922
rect 1972 4868 1996 4870
rect 2052 4868 2076 4870
rect 2132 4868 2156 4870
rect 2212 4868 2236 4870
rect 1916 4859 2292 4868
rect 2656 4380 3032 4389
rect 2712 4378 2736 4380
rect 2792 4378 2816 4380
rect 2872 4378 2896 4380
rect 2952 4378 2976 4380
rect 2712 4326 2722 4378
rect 2966 4326 2976 4378
rect 2712 4324 2736 4326
rect 2792 4324 2816 4326
rect 2872 4324 2896 4326
rect 2952 4324 2976 4326
rect 2656 4315 3032 4324
rect 3436 4146 3464 10628
rect 3528 10198 3556 11494
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3620 9518 3648 11154
rect 3700 11076 3752 11082
rect 3700 11018 3752 11024
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3712 9364 3740 11018
rect 3528 9336 3740 9364
rect 3528 8974 3556 9336
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 3528 8378 3556 8910
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3620 8566 3648 8774
rect 3608 8560 3660 8566
rect 3608 8502 3660 8508
rect 3700 8560 3752 8566
rect 3700 8502 3752 8508
rect 3528 8350 3648 8378
rect 3620 8294 3648 8350
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3528 8090 3556 8230
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3620 7562 3648 8026
rect 3528 7534 3648 7562
rect 3528 6225 3556 7534
rect 3608 7472 3660 7478
rect 3608 7414 3660 7420
rect 3514 6216 3570 6225
rect 3514 6151 3570 6160
rect 3620 5681 3648 7414
rect 3606 5672 3662 5681
rect 3516 5636 3568 5642
rect 3606 5607 3662 5616
rect 3516 5578 3568 5584
rect 3528 5166 3556 5578
rect 3712 5370 3740 8502
rect 3804 7886 3832 12815
rect 4264 12434 4292 15399
rect 4448 15162 4476 17138
rect 4540 15910 4568 17206
rect 4816 17202 4844 19314
rect 4908 18222 4936 20810
rect 5356 20800 5408 20806
rect 5356 20742 5408 20748
rect 5368 20466 5396 20742
rect 5552 20482 5580 20946
rect 5460 20466 5580 20482
rect 5356 20460 5408 20466
rect 5356 20402 5408 20408
rect 5448 20460 5580 20466
rect 5500 20454 5580 20460
rect 5448 20402 5500 20408
rect 5644 20058 5672 21490
rect 6552 21480 6604 21486
rect 6552 21422 6604 21428
rect 6564 21010 6592 21422
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 6552 21004 6604 21010
rect 6552 20946 6604 20952
rect 5632 20052 5684 20058
rect 5632 19994 5684 20000
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 5276 19514 5304 19654
rect 5264 19508 5316 19514
rect 5264 19450 5316 19456
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 5092 18970 5120 19314
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 5920 18766 5948 19110
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 5908 18760 5960 18766
rect 5908 18702 5960 18708
rect 5368 18426 5396 18702
rect 5540 18692 5592 18698
rect 5540 18634 5592 18640
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4620 17060 4672 17066
rect 4620 17002 4672 17008
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4540 15502 4568 15846
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4632 15094 4660 17002
rect 4908 16182 4936 18022
rect 5354 17776 5410 17785
rect 5354 17711 5410 17720
rect 5368 17678 5396 17711
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 4896 16176 4948 16182
rect 4896 16118 4948 16124
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4724 15706 4752 15982
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4816 15609 4844 15642
rect 4802 15600 4858 15609
rect 4802 15535 4858 15544
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4620 15088 4672 15094
rect 4620 15030 4672 15036
rect 4724 14346 4752 15370
rect 5092 15162 5120 17138
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 5184 16658 5212 16934
rect 5172 16652 5224 16658
rect 5172 16594 5224 16600
rect 5460 16454 5488 18362
rect 5552 18290 5580 18634
rect 6196 18290 6224 20946
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6644 20460 6696 20466
rect 6644 20402 6696 20408
rect 6276 20324 6328 20330
rect 6276 20266 6328 20272
rect 6288 19786 6316 20266
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 6380 19786 6408 20198
rect 6564 20058 6592 20198
rect 6552 20052 6604 20058
rect 6552 19994 6604 20000
rect 6276 19780 6328 19786
rect 6276 19722 6328 19728
rect 6368 19780 6420 19786
rect 6368 19722 6420 19728
rect 6288 18358 6316 19722
rect 6276 18352 6328 18358
rect 6276 18294 6328 18300
rect 5540 18284 5592 18290
rect 5540 18226 5592 18232
rect 6092 18284 6144 18290
rect 6092 18226 6144 18232
rect 6184 18284 6236 18290
rect 6184 18226 6236 18232
rect 5908 16992 5960 16998
rect 5828 16940 5908 16946
rect 5828 16934 5960 16940
rect 5828 16918 5948 16934
rect 5828 16590 5856 16918
rect 6104 16794 6132 18226
rect 6196 16794 6224 18226
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5354 16008 5410 16017
rect 5410 15966 5488 15994
rect 5354 15943 5410 15952
rect 5460 15638 5488 15966
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 6104 15162 6132 16730
rect 6288 16590 6316 18022
rect 6552 17604 6604 17610
rect 6552 17546 6604 17552
rect 6564 17338 6592 17546
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 6368 17264 6420 17270
rect 6368 17206 6420 17212
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 6380 15910 6408 17206
rect 6460 16992 6512 16998
rect 6460 16934 6512 16940
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 5080 15156 5132 15162
rect 5080 15098 5132 15104
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 5092 14550 5120 15098
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 5080 14544 5132 14550
rect 5080 14486 5132 14492
rect 4436 14340 4488 14346
rect 4436 14282 4488 14288
rect 4712 14340 4764 14346
rect 4712 14282 4764 14288
rect 4448 13938 4476 14282
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 4356 13138 4384 13194
rect 4356 13110 4660 13138
rect 4632 12714 4660 13110
rect 4816 12986 4844 13806
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 4264 12406 4384 12434
rect 4356 12306 4384 12406
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 3976 12164 4028 12170
rect 3976 12106 4028 12112
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3896 10198 3924 10610
rect 3884 10192 3936 10198
rect 3884 10134 3936 10140
rect 3988 9058 4016 12106
rect 4172 9586 4200 12106
rect 4344 11620 4396 11626
rect 4344 11562 4396 11568
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 3896 9030 4016 9058
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3790 7712 3846 7721
rect 3790 7647 3846 7656
rect 3804 7546 3832 7647
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3804 6497 3832 6734
rect 3790 6488 3846 6497
rect 3790 6423 3846 6432
rect 3804 5846 3832 6423
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3804 5370 3832 5782
rect 3896 5574 3924 9030
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3988 8566 4016 8910
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 4080 7154 4108 8910
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 3988 7126 4108 7154
rect 3988 6848 4016 7126
rect 4172 7002 4200 7414
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4264 6866 4292 10542
rect 4356 10130 4384 11562
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4356 7818 4384 8842
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4342 7304 4398 7313
rect 4448 7274 4476 11086
rect 4528 11076 4580 11082
rect 4528 11018 4580 11024
rect 4540 9994 4568 11018
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4724 9926 4752 12854
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4908 12170 4936 12786
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4816 10713 4844 11018
rect 4802 10704 4858 10713
rect 4802 10639 4858 10648
rect 5092 10470 5120 13874
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5368 12986 5396 13126
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5460 11150 5488 13126
rect 5644 11354 5672 13874
rect 6380 13802 6408 14758
rect 6472 14414 6500 16934
rect 6656 16114 6684 20402
rect 6748 18970 6776 20878
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6840 18834 6868 21830
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 7012 20800 7064 20806
rect 7012 20742 7064 20748
rect 6828 18828 6880 18834
rect 6828 18770 6880 18776
rect 6932 18766 6960 20742
rect 7024 19446 7052 20742
rect 7576 19514 7604 24142
rect 8656 23964 9032 23973
rect 8712 23962 8736 23964
rect 8792 23962 8816 23964
rect 8872 23962 8896 23964
rect 8952 23962 8976 23964
rect 8712 23910 8722 23962
rect 8966 23910 8976 23962
rect 8712 23908 8736 23910
rect 8792 23908 8816 23910
rect 8872 23908 8896 23910
rect 8952 23908 8976 23910
rect 8656 23899 9032 23908
rect 7916 23420 8292 23429
rect 7972 23418 7996 23420
rect 8052 23418 8076 23420
rect 8132 23418 8156 23420
rect 8212 23418 8236 23420
rect 7972 23366 7982 23418
rect 8226 23366 8236 23418
rect 7972 23364 7996 23366
rect 8052 23364 8076 23366
rect 8132 23364 8156 23366
rect 8212 23364 8236 23366
rect 7916 23355 8292 23364
rect 8656 22876 9032 22885
rect 8712 22874 8736 22876
rect 8792 22874 8816 22876
rect 8872 22874 8896 22876
rect 8952 22874 8976 22876
rect 8712 22822 8722 22874
rect 8966 22822 8976 22874
rect 8712 22820 8736 22822
rect 8792 22820 8816 22822
rect 8872 22820 8896 22822
rect 8952 22820 8976 22822
rect 8656 22811 9032 22820
rect 7916 22332 8292 22341
rect 7972 22330 7996 22332
rect 8052 22330 8076 22332
rect 8132 22330 8156 22332
rect 8212 22330 8236 22332
rect 7972 22278 7982 22330
rect 8226 22278 8236 22330
rect 7972 22276 7996 22278
rect 8052 22276 8076 22278
rect 8132 22276 8156 22278
rect 8212 22276 8236 22278
rect 7916 22267 8292 22276
rect 7840 21956 7892 21962
rect 7840 21898 7892 21904
rect 7656 21480 7708 21486
rect 7656 21422 7708 21428
rect 7668 20262 7696 21422
rect 7748 21344 7800 21350
rect 7748 21286 7800 21292
rect 7760 20466 7788 21286
rect 7852 20942 7880 21898
rect 8576 21888 8628 21894
rect 8576 21830 8628 21836
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 7916 21244 8292 21253
rect 7972 21242 7996 21244
rect 8052 21242 8076 21244
rect 8132 21242 8156 21244
rect 8212 21242 8236 21244
rect 7972 21190 7982 21242
rect 8226 21190 8236 21242
rect 7972 21188 7996 21190
rect 8052 21188 8076 21190
rect 8132 21188 8156 21190
rect 8212 21188 8236 21190
rect 7916 21179 8292 21188
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 7840 20800 7892 20806
rect 7840 20742 7892 20748
rect 8300 20800 8352 20806
rect 8300 20742 8352 20748
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 7852 19786 7880 20742
rect 8312 20602 8340 20742
rect 8300 20596 8352 20602
rect 8300 20538 8352 20544
rect 7916 20156 8292 20165
rect 7972 20154 7996 20156
rect 8052 20154 8076 20156
rect 8132 20154 8156 20156
rect 8212 20154 8236 20156
rect 7972 20102 7982 20154
rect 8226 20102 8236 20154
rect 7972 20100 7996 20102
rect 8052 20100 8076 20102
rect 8132 20100 8156 20102
rect 8212 20100 8236 20102
rect 7916 20091 8292 20100
rect 7840 19780 7892 19786
rect 7840 19722 7892 19728
rect 8300 19780 8352 19786
rect 8300 19722 8352 19728
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 7012 19440 7064 19446
rect 7012 19382 7064 19388
rect 8312 19394 8340 19722
rect 8404 19514 8432 20742
rect 8496 19938 8524 21286
rect 8588 20466 8616 21830
rect 8656 21788 9032 21797
rect 8712 21786 8736 21788
rect 8792 21786 8816 21788
rect 8872 21786 8896 21788
rect 8952 21786 8976 21788
rect 8712 21734 8722 21786
rect 8966 21734 8976 21786
rect 8712 21732 8736 21734
rect 8792 21732 8816 21734
rect 8872 21732 8896 21734
rect 8952 21732 8976 21734
rect 8656 21723 9032 21732
rect 9496 21480 9548 21486
rect 9496 21422 9548 21428
rect 9312 21344 9364 21350
rect 9312 21286 9364 21292
rect 9404 21344 9456 21350
rect 9404 21286 9456 21292
rect 9220 20868 9272 20874
rect 9220 20810 9272 20816
rect 9128 20800 9180 20806
rect 9128 20742 9180 20748
rect 8656 20700 9032 20709
rect 8712 20698 8736 20700
rect 8792 20698 8816 20700
rect 8872 20698 8896 20700
rect 8952 20698 8976 20700
rect 8712 20646 8722 20698
rect 8966 20646 8976 20698
rect 8712 20644 8736 20646
rect 8792 20644 8816 20646
rect 8872 20644 8896 20646
rect 8952 20644 8976 20646
rect 8656 20635 9032 20644
rect 8668 20596 8720 20602
rect 8668 20538 8720 20544
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 8496 19910 8616 19938
rect 8588 19854 8616 19910
rect 8680 19854 8708 20538
rect 9140 19922 9168 20742
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 8484 19848 8536 19854
rect 8484 19790 8536 19796
rect 8576 19848 8628 19854
rect 8576 19790 8628 19796
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 8392 19508 8444 19514
rect 8392 19450 8444 19456
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6748 17338 6776 18226
rect 7024 17746 7052 19382
rect 8312 19378 8432 19394
rect 8312 19372 8444 19378
rect 8312 19366 8392 19372
rect 8392 19314 8444 19320
rect 7916 19068 8292 19077
rect 7972 19066 7996 19068
rect 8052 19066 8076 19068
rect 8132 19066 8156 19068
rect 8212 19066 8236 19068
rect 7972 19014 7982 19066
rect 8226 19014 8236 19066
rect 7972 19012 7996 19014
rect 8052 19012 8076 19014
rect 8132 19012 8156 19014
rect 8212 19012 8236 19014
rect 7916 19003 8292 19012
rect 8496 18766 8524 19790
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7484 17882 7512 18226
rect 7840 18148 7892 18154
rect 7840 18090 7892 18096
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7012 17740 7064 17746
rect 7012 17682 7064 17688
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6736 17332 6788 17338
rect 6736 17274 6788 17280
rect 6840 16794 6868 17478
rect 6932 17338 6960 17478
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6840 14074 6868 15846
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 5816 13252 5868 13258
rect 5816 13194 5868 13200
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5828 11218 5856 13194
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6196 12434 6224 12582
rect 5920 12406 6224 12434
rect 5920 11762 5948 12406
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5552 10810 5580 11086
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 6000 9988 6052 9994
rect 6000 9930 6052 9936
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4724 9586 4752 9862
rect 5552 9586 5580 9930
rect 6012 9722 6040 9930
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4342 7239 4398 7248
rect 4436 7268 4488 7274
rect 4252 6860 4304 6866
rect 3988 6820 4108 6848
rect 3974 6624 4030 6633
rect 3974 6559 4030 6568
rect 3988 5953 4016 6559
rect 3974 5944 4030 5953
rect 4080 5914 4108 6820
rect 4252 6802 4304 6808
rect 4356 6322 4384 7239
rect 4436 7210 4488 7216
rect 4540 6905 4568 8230
rect 4632 7206 4660 9522
rect 4724 8974 4752 9522
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4526 6896 4582 6905
rect 4526 6831 4582 6840
rect 4540 6390 4568 6831
rect 4632 6769 4660 6938
rect 4618 6760 4674 6769
rect 4618 6695 4674 6704
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4724 6322 4752 8910
rect 4816 7721 4844 9454
rect 5092 9178 5120 9522
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4908 7886 4936 8230
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4988 7812 5040 7818
rect 4988 7754 5040 7760
rect 4802 7712 4858 7721
rect 4802 7647 4858 7656
rect 5000 7410 5028 7754
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4344 6180 4396 6186
rect 4344 6122 4396 6128
rect 4356 6066 4384 6122
rect 4264 6038 4384 6066
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4264 5914 4292 6038
rect 3974 5879 4030 5888
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 3976 5704 4028 5710
rect 4028 5664 4108 5692
rect 3976 5646 4028 5652
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3988 5234 4016 5510
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 4080 4690 4108 5664
rect 4448 5234 4476 6054
rect 4632 5642 4660 6258
rect 4724 5642 4752 6258
rect 4620 5636 4672 5642
rect 4620 5578 4672 5584
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4632 5370 4660 5578
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4908 5234 4936 7346
rect 5092 5574 5120 8910
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 5184 8090 5212 8502
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5460 7970 5488 8774
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5276 7942 5488 7970
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 1916 3836 2292 3845
rect 1972 3834 1996 3836
rect 2052 3834 2076 3836
rect 2132 3834 2156 3836
rect 2212 3834 2236 3836
rect 1972 3782 1982 3834
rect 2226 3782 2236 3834
rect 1972 3780 1996 3782
rect 2052 3780 2076 3782
rect 2132 3780 2156 3782
rect 2212 3780 2236 3782
rect 1916 3771 2292 3780
rect 2656 3292 3032 3301
rect 2712 3290 2736 3292
rect 2792 3290 2816 3292
rect 2872 3290 2896 3292
rect 2952 3290 2976 3292
rect 2712 3238 2722 3290
rect 2966 3238 2976 3290
rect 2712 3236 2736 3238
rect 2792 3236 2816 3238
rect 2872 3236 2896 3238
rect 2952 3236 2976 3238
rect 2656 3227 3032 3236
rect 5276 2774 5304 7942
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5368 7041 5396 7754
rect 5460 7177 5488 7822
rect 5552 7206 5580 8434
rect 5644 7886 5672 8842
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5920 7410 5948 8230
rect 6104 7546 6132 11698
rect 6288 10010 6316 12038
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6380 10266 6408 11630
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6288 9982 6408 10010
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5540 7200 5592 7206
rect 5446 7168 5502 7177
rect 5540 7142 5592 7148
rect 5446 7103 5502 7112
rect 5354 7032 5410 7041
rect 5354 6967 5410 6976
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5828 4826 5856 6734
rect 6196 6458 6224 8366
rect 6288 7410 6316 9862
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 6012 4622 6040 5170
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6012 4282 6040 4558
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 1916 2748 2292 2757
rect 1972 2746 1996 2748
rect 2052 2746 2076 2748
rect 2132 2746 2156 2748
rect 2212 2746 2236 2748
rect 5276 2746 5488 2774
rect 1972 2694 1982 2746
rect 2226 2694 2236 2746
rect 1972 2692 1996 2694
rect 2052 2692 2076 2694
rect 2132 2692 2156 2694
rect 2212 2692 2236 2694
rect 1916 2683 2292 2692
rect 5460 2446 5488 2746
rect 6288 2582 6316 6598
rect 6380 3058 6408 9982
rect 6472 9625 6500 10610
rect 6458 9616 6514 9625
rect 6458 9551 6514 9560
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6472 5817 6500 8230
rect 6564 7478 6592 8774
rect 6552 7472 6604 7478
rect 6552 7414 6604 7420
rect 6656 6458 6684 13262
rect 6932 12968 6960 17274
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7012 17060 7064 17066
rect 7012 17002 7064 17008
rect 7024 16114 7052 17002
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 7012 15972 7064 15978
rect 7012 15914 7064 15920
rect 7024 13462 7052 15914
rect 7116 15162 7144 17070
rect 7484 15706 7512 17818
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 6748 12940 6960 12968
rect 6748 12782 6776 12940
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6748 6361 6776 9658
rect 6840 9654 6868 12786
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6840 6662 6868 7278
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6932 6497 6960 10406
rect 7024 6769 7052 13398
rect 7116 9450 7144 14214
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7208 12850 7236 13126
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7196 12164 7248 12170
rect 7196 12106 7248 12112
rect 7208 10266 7236 12106
rect 7300 10742 7328 14214
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7668 12714 7696 12786
rect 7656 12708 7708 12714
rect 7656 12650 7708 12656
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7484 12102 7512 12582
rect 7576 12434 7604 12582
rect 7656 12436 7708 12442
rect 7576 12406 7656 12434
rect 7656 12378 7708 12384
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7668 11150 7696 11494
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7288 10736 7340 10742
rect 7288 10678 7340 10684
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 7116 7993 7144 9386
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7208 8566 7236 9318
rect 7196 8560 7248 8566
rect 7196 8502 7248 8508
rect 7102 7984 7158 7993
rect 7102 7919 7158 7928
rect 7392 7546 7420 11086
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7484 10742 7512 10950
rect 7472 10736 7524 10742
rect 7472 10678 7524 10684
rect 7760 10198 7788 16390
rect 7852 16114 7880 18090
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 7916 17980 8292 17989
rect 7972 17978 7996 17980
rect 8052 17978 8076 17980
rect 8132 17978 8156 17980
rect 8212 17978 8236 17980
rect 7972 17926 7982 17978
rect 8226 17926 8236 17978
rect 7972 17924 7996 17926
rect 8052 17924 8076 17926
rect 8132 17924 8156 17926
rect 8212 17924 8236 17926
rect 7916 17915 8292 17924
rect 7916 16892 8292 16901
rect 7972 16890 7996 16892
rect 8052 16890 8076 16892
rect 8132 16890 8156 16892
rect 8212 16890 8236 16892
rect 7972 16838 7982 16890
rect 8226 16838 8236 16890
rect 7972 16836 7996 16838
rect 8052 16836 8076 16838
rect 8132 16836 8156 16838
rect 8212 16836 8236 16838
rect 7916 16827 8292 16836
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 8312 16017 8340 16390
rect 8298 16008 8354 16017
rect 8298 15943 8354 15952
rect 7916 15804 8292 15813
rect 7972 15802 7996 15804
rect 8052 15802 8076 15804
rect 8132 15802 8156 15804
rect 8212 15802 8236 15804
rect 7972 15750 7982 15802
rect 8226 15750 8236 15802
rect 7972 15748 7996 15750
rect 8052 15748 8076 15750
rect 8132 15748 8156 15750
rect 8212 15748 8236 15750
rect 7916 15739 8292 15748
rect 8404 15434 8432 18022
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8392 15428 8444 15434
rect 8392 15370 8444 15376
rect 8496 15162 8524 17546
rect 8588 15706 8616 19654
rect 8656 19612 9032 19621
rect 8712 19610 8736 19612
rect 8792 19610 8816 19612
rect 8872 19610 8896 19612
rect 8952 19610 8976 19612
rect 8712 19558 8722 19610
rect 8966 19558 8976 19610
rect 8712 19556 8736 19558
rect 8792 19556 8816 19558
rect 8872 19556 8896 19558
rect 8952 19556 8976 19558
rect 8656 19547 9032 19556
rect 9232 19378 9260 20810
rect 9324 20534 9352 21286
rect 9416 20806 9444 21286
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 9312 20528 9364 20534
rect 9312 20470 9364 20476
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9220 19372 9272 19378
rect 9220 19314 9272 19320
rect 8656 18524 9032 18533
rect 8712 18522 8736 18524
rect 8792 18522 8816 18524
rect 8872 18522 8896 18524
rect 8952 18522 8976 18524
rect 8712 18470 8722 18522
rect 8966 18470 8976 18522
rect 8712 18468 8736 18470
rect 8792 18468 8816 18470
rect 8872 18468 8896 18470
rect 8952 18468 8976 18470
rect 8656 18459 9032 18468
rect 9324 18426 9352 19790
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 8656 17436 9032 17445
rect 8712 17434 8736 17436
rect 8792 17434 8816 17436
rect 8872 17434 8896 17436
rect 8952 17434 8976 17436
rect 8712 17382 8722 17434
rect 8966 17382 8976 17434
rect 8712 17380 8736 17382
rect 8792 17380 8816 17382
rect 8872 17380 8896 17382
rect 8952 17380 8976 17382
rect 8656 17371 9032 17380
rect 8666 17096 8722 17105
rect 8666 17031 8722 17040
rect 8680 16522 8708 17031
rect 9036 16720 9088 16726
rect 9034 16688 9036 16697
rect 9088 16688 9090 16697
rect 9034 16623 9090 16632
rect 8668 16516 8720 16522
rect 8668 16458 8720 16464
rect 8656 16348 9032 16357
rect 8712 16346 8736 16348
rect 8792 16346 8816 16348
rect 8872 16346 8896 16348
rect 8952 16346 8976 16348
rect 8712 16294 8722 16346
rect 8966 16294 8976 16346
rect 8712 16292 8736 16294
rect 8792 16292 8816 16294
rect 8872 16292 8896 16294
rect 8952 16292 8976 16294
rect 8656 16283 9032 16292
rect 9140 16153 9168 17614
rect 9416 17338 9444 20742
rect 9508 19990 9536 21422
rect 9600 20618 9628 24142
rect 10324 22160 10376 22166
rect 10324 22102 10376 22108
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 9600 20590 9720 20618
rect 9588 20460 9640 20466
rect 9588 20402 9640 20408
rect 9600 19990 9628 20402
rect 9496 19984 9548 19990
rect 9496 19926 9548 19932
rect 9588 19984 9640 19990
rect 9588 19926 9640 19932
rect 9496 19848 9548 19854
rect 9692 19836 9720 20590
rect 9496 19790 9548 19796
rect 9600 19808 9720 19836
rect 9508 19514 9536 19790
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9600 18902 9628 19808
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9588 18896 9640 18902
rect 9588 18838 9640 18844
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9126 16144 9182 16153
rect 9126 16079 9182 16088
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8656 15260 9032 15269
rect 8712 15258 8736 15260
rect 8792 15258 8816 15260
rect 8872 15258 8896 15260
rect 8952 15258 8976 15260
rect 8712 15206 8722 15258
rect 8966 15206 8976 15258
rect 8712 15204 8736 15206
rect 8792 15204 8816 15206
rect 8872 15204 8896 15206
rect 8952 15204 8976 15206
rect 8656 15195 9032 15204
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 7916 14716 8292 14725
rect 7972 14714 7996 14716
rect 8052 14714 8076 14716
rect 8132 14714 8156 14716
rect 8212 14714 8236 14716
rect 7972 14662 7982 14714
rect 8226 14662 8236 14714
rect 7972 14660 7996 14662
rect 8052 14660 8076 14662
rect 8132 14660 8156 14662
rect 8212 14660 8236 14662
rect 7916 14651 8292 14660
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 7916 13628 8292 13637
rect 7972 13626 7996 13628
rect 8052 13626 8076 13628
rect 8132 13626 8156 13628
rect 8212 13626 8236 13628
rect 7972 13574 7982 13626
rect 8226 13574 8236 13626
rect 7972 13572 7996 13574
rect 8052 13572 8076 13574
rect 8132 13572 8156 13574
rect 8212 13572 8236 13574
rect 7916 13563 8292 13572
rect 8404 13258 8432 13806
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8496 12968 8524 15098
rect 8656 14172 9032 14181
rect 8712 14170 8736 14172
rect 8792 14170 8816 14172
rect 8872 14170 8896 14172
rect 8952 14170 8976 14172
rect 8712 14118 8722 14170
rect 8966 14118 8976 14170
rect 8712 14116 8736 14118
rect 8792 14116 8816 14118
rect 8872 14116 8896 14118
rect 8952 14116 8976 14118
rect 8656 14107 9032 14116
rect 9140 14056 9168 16079
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 9232 14634 9260 15302
rect 9232 14606 9352 14634
rect 9048 14028 9168 14056
rect 9048 13258 9076 14028
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 8656 13084 9032 13093
rect 8712 13082 8736 13084
rect 8792 13082 8816 13084
rect 8872 13082 8896 13084
rect 8952 13082 8976 13084
rect 8712 13030 8722 13082
rect 8966 13030 8976 13082
rect 8712 13028 8736 13030
rect 8792 13028 8816 13030
rect 8872 13028 8896 13030
rect 8952 13028 8976 13030
rect 8656 13019 9032 13028
rect 8496 12940 8708 12968
rect 8390 12880 8446 12889
rect 8390 12815 8392 12824
rect 8444 12815 8446 12824
rect 8392 12786 8444 12792
rect 7916 12540 8292 12549
rect 7972 12538 7996 12540
rect 8052 12538 8076 12540
rect 8132 12538 8156 12540
rect 8212 12538 8236 12540
rect 7972 12486 7982 12538
rect 8226 12486 8236 12538
rect 7972 12484 7996 12486
rect 8052 12484 8076 12486
rect 8132 12484 8156 12486
rect 8212 12484 8236 12486
rect 7916 12475 8292 12484
rect 8680 12434 8708 12940
rect 8680 12406 8984 12434
rect 8956 12238 8984 12406
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8392 12164 8444 12170
rect 8392 12106 8444 12112
rect 7916 11452 8292 11461
rect 7972 11450 7996 11452
rect 8052 11450 8076 11452
rect 8132 11450 8156 11452
rect 8212 11450 8236 11452
rect 7972 11398 7982 11450
rect 8226 11398 8236 11450
rect 7972 11396 7996 11398
rect 8052 11396 8076 11398
rect 8132 11396 8156 11398
rect 8212 11396 8236 11398
rect 7916 11387 8292 11396
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7852 10130 7880 10610
rect 7916 10364 8292 10373
rect 7972 10362 7996 10364
rect 8052 10362 8076 10364
rect 8132 10362 8156 10364
rect 8212 10362 8236 10364
rect 7972 10310 7982 10362
rect 8226 10310 8236 10362
rect 7972 10308 7996 10310
rect 8052 10308 8076 10310
rect 8132 10308 8156 10310
rect 8212 10308 8236 10310
rect 7916 10299 8292 10308
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7852 8566 7880 10066
rect 7916 9276 8292 9285
rect 7972 9274 7996 9276
rect 8052 9274 8076 9276
rect 8132 9274 8156 9276
rect 8212 9274 8236 9276
rect 7972 9222 7982 9274
rect 8226 9222 8236 9274
rect 7972 9220 7996 9222
rect 8052 9220 8076 9222
rect 8132 9220 8156 9222
rect 8212 9220 8236 9222
rect 7916 9211 8292 9220
rect 8404 9178 8432 12106
rect 8656 11996 9032 12005
rect 8712 11994 8736 11996
rect 8792 11994 8816 11996
rect 8872 11994 8896 11996
rect 8952 11994 8976 11996
rect 8712 11942 8722 11994
rect 8966 11942 8976 11994
rect 8712 11940 8736 11942
rect 8792 11940 8816 11942
rect 8872 11940 8896 11942
rect 8952 11940 8976 11942
rect 8656 11931 9032 11940
rect 9140 11558 9168 13874
rect 9324 13274 9352 14606
rect 9232 13246 9352 13274
rect 9232 12170 9260 13246
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9220 12164 9272 12170
rect 9220 12106 9272 12112
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 8496 10742 8524 11494
rect 9324 11098 9352 13126
rect 9416 12753 9444 16458
rect 9508 15978 9536 18634
rect 9692 17746 9720 19654
rect 9784 19174 9812 21422
rect 9968 20398 9996 21966
rect 9956 20392 10008 20398
rect 9956 20334 10008 20340
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 9876 18970 9904 19790
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9968 18306 9996 20334
rect 10060 18970 10088 22034
rect 10336 21690 10364 22102
rect 10508 21956 10560 21962
rect 10508 21898 10560 21904
rect 10600 21956 10652 21962
rect 10600 21898 10652 21904
rect 10520 21690 10548 21898
rect 10324 21684 10376 21690
rect 10324 21626 10376 21632
rect 10508 21684 10560 21690
rect 10508 21626 10560 21632
rect 10508 21548 10560 21554
rect 10508 21490 10560 21496
rect 10416 21480 10468 21486
rect 10416 21422 10468 21428
rect 10428 20602 10456 21422
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 10060 18426 10088 18566
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 9876 18278 9996 18306
rect 9876 18222 9904 18278
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9876 16454 9904 18158
rect 10152 17785 10180 19314
rect 10520 18766 10548 21490
rect 10612 20874 10640 21898
rect 10600 20868 10652 20874
rect 10600 20810 10652 20816
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10508 18760 10560 18766
rect 10508 18702 10560 18708
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10612 17882 10640 18226
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10138 17776 10194 17785
rect 10138 17711 10194 17720
rect 10704 17610 10732 19314
rect 10796 19310 10824 24142
rect 10968 22432 11020 22438
rect 10968 22374 11020 22380
rect 10980 22094 11008 22374
rect 10888 22066 11008 22094
rect 10888 19786 10916 22066
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 10968 21956 11020 21962
rect 10968 21898 11020 21904
rect 10980 21146 11008 21898
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 12072 21888 12124 21894
rect 12072 21830 12124 21836
rect 11072 21622 11100 21830
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 11060 21616 11112 21622
rect 11060 21558 11112 21564
rect 10968 21140 11020 21146
rect 10968 21082 11020 21088
rect 11072 20806 11100 21558
rect 11612 21548 11664 21554
rect 11532 21508 11612 21536
rect 11152 21344 11204 21350
rect 11152 21286 11204 21292
rect 11244 21344 11296 21350
rect 11244 21286 11296 21292
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 10876 19780 10928 19786
rect 10876 19722 10928 19728
rect 11072 19310 11100 20742
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10692 17604 10744 17610
rect 10692 17546 10744 17552
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9508 14278 9536 15914
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9402 12744 9458 12753
rect 9402 12679 9458 12688
rect 9404 12640 9456 12646
rect 9402 12608 9404 12617
rect 9456 12608 9458 12617
rect 9402 12543 9458 12552
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 9232 11082 9352 11098
rect 9128 11076 9180 11082
rect 9128 11018 9180 11024
rect 9220 11076 9352 11082
rect 9272 11070 9352 11076
rect 9220 11018 9272 11024
rect 8656 10908 9032 10917
rect 8712 10906 8736 10908
rect 8792 10906 8816 10908
rect 8872 10906 8896 10908
rect 8952 10906 8976 10908
rect 8712 10854 8722 10906
rect 8966 10854 8976 10906
rect 8712 10852 8736 10854
rect 8792 10852 8816 10854
rect 8872 10852 8896 10854
rect 8952 10852 8976 10854
rect 8656 10843 9032 10852
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8496 8974 8524 9862
rect 8656 9820 9032 9829
rect 8712 9818 8736 9820
rect 8792 9818 8816 9820
rect 8872 9818 8896 9820
rect 8952 9818 8976 9820
rect 8712 9766 8722 9818
rect 8966 9766 8976 9818
rect 8712 9764 8736 9766
rect 8792 9764 8816 9766
rect 8872 9764 8896 9766
rect 8952 9764 8976 9766
rect 8656 9755 9032 9764
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7916 8188 8292 8197
rect 7972 8186 7996 8188
rect 8052 8186 8076 8188
rect 8132 8186 8156 8188
rect 8212 8186 8236 8188
rect 7972 8134 7982 8186
rect 8226 8134 8236 8186
rect 7972 8132 7996 8134
rect 8052 8132 8076 8134
rect 8132 8132 8156 8134
rect 8212 8132 8236 8134
rect 7916 8123 8292 8132
rect 7472 7880 7524 7886
rect 8588 7857 8616 8842
rect 8656 8732 9032 8741
rect 8712 8730 8736 8732
rect 8792 8730 8816 8732
rect 8872 8730 8896 8732
rect 8952 8730 8976 8732
rect 8712 8678 8722 8730
rect 8966 8678 8976 8730
rect 8712 8676 8736 8678
rect 8792 8676 8816 8678
rect 8872 8676 8896 8678
rect 8952 8676 8976 8678
rect 8656 8667 9032 8676
rect 8944 8424 8996 8430
rect 8944 8366 8996 8372
rect 8956 8090 8984 8366
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 7472 7822 7524 7828
rect 8574 7848 8630 7857
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7288 6792 7340 6798
rect 7010 6760 7066 6769
rect 7288 6734 7340 6740
rect 7010 6695 7066 6704
rect 6918 6488 6974 6497
rect 7024 6458 7052 6695
rect 6918 6423 6920 6432
rect 6972 6423 6974 6432
rect 7012 6452 7064 6458
rect 6920 6394 6972 6400
rect 7012 6394 7064 6400
rect 6734 6352 6790 6361
rect 6734 6287 6790 6296
rect 7104 6316 7156 6322
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6458 5808 6514 5817
rect 6458 5743 6514 5752
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 6472 5302 6500 5578
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6564 4146 6592 6190
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6656 4622 6684 6054
rect 6748 4622 6776 6287
rect 7104 6258 7156 6264
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6840 4162 6868 5510
rect 7116 4622 7144 6258
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 6840 4146 6960 4162
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6552 4140 6604 4146
rect 6840 4140 6972 4146
rect 6840 4134 6920 4140
rect 6552 4082 6604 4088
rect 6920 4082 6972 4088
rect 6472 3534 6500 4082
rect 7208 3738 7236 5646
rect 7300 5370 7328 6734
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7392 5250 7420 5510
rect 7300 5222 7420 5250
rect 7300 3942 7328 5222
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7392 4826 7420 5102
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7484 3670 7512 7822
rect 8574 7783 8630 7792
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7852 7546 7880 7686
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 8128 7500 8340 7528
rect 8128 7206 8156 7500
rect 8312 7410 8340 7500
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8220 7206 8248 7346
rect 8404 7342 8432 7414
rect 8392 7336 8444 7342
rect 8444 7284 8524 7290
rect 8392 7278 8524 7284
rect 8404 7262 8524 7278
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 7916 7100 8292 7109
rect 7972 7098 7996 7100
rect 8052 7098 8076 7100
rect 8132 7098 8156 7100
rect 8212 7098 8236 7100
rect 7972 7046 7982 7098
rect 8226 7046 8236 7098
rect 7972 7044 7996 7046
rect 8052 7044 8076 7046
rect 8132 7044 8156 7046
rect 8212 7044 8236 7046
rect 7916 7035 8292 7044
rect 8404 7002 8432 7142
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 7656 6724 7708 6730
rect 7656 6666 7708 6672
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7576 4826 7604 6258
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7668 4622 7696 6666
rect 8312 6225 8340 6870
rect 8496 6866 8524 7262
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8298 6216 8354 6225
rect 8298 6151 8354 6160
rect 7916 6012 8292 6021
rect 7972 6010 7996 6012
rect 8052 6010 8076 6012
rect 8132 6010 8156 6012
rect 8212 6010 8236 6012
rect 7972 5958 7982 6010
rect 8226 5958 8236 6010
rect 7972 5956 7996 5958
rect 8052 5956 8076 5958
rect 8132 5956 8156 5958
rect 8212 5956 8236 5958
rect 7916 5947 8292 5956
rect 8496 5710 8524 6598
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7760 4622 7788 4966
rect 7916 4924 8292 4933
rect 7972 4922 7996 4924
rect 8052 4922 8076 4924
rect 8132 4922 8156 4924
rect 8212 4922 8236 4924
rect 7972 4870 7982 4922
rect 8226 4870 8236 4922
rect 7972 4868 7996 4870
rect 8052 4868 8076 4870
rect 8132 4868 8156 4870
rect 8212 4868 8236 4870
rect 7916 4859 8292 4868
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8128 4282 8156 4422
rect 8312 4282 8340 4558
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 7916 3836 8292 3845
rect 7972 3834 7996 3836
rect 8052 3834 8076 3836
rect 8132 3834 8156 3836
rect 8212 3834 8236 3836
rect 7972 3782 7982 3834
rect 8226 3782 8236 3834
rect 7972 3780 7996 3782
rect 8052 3780 8076 3782
rect 8132 3780 8156 3782
rect 8212 3780 8236 3782
rect 7916 3771 8292 3780
rect 8404 3738 8432 5646
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 8496 3534 8524 4490
rect 8588 4146 8616 7783
rect 8656 7644 9032 7653
rect 8712 7642 8736 7644
rect 8792 7642 8816 7644
rect 8872 7642 8896 7644
rect 8952 7642 8976 7644
rect 8712 7590 8722 7642
rect 8966 7590 8976 7642
rect 8712 7588 8736 7590
rect 8792 7588 8816 7590
rect 8872 7588 8896 7590
rect 8952 7588 8976 7590
rect 8656 7579 9032 7588
rect 8656 6556 9032 6565
rect 8712 6554 8736 6556
rect 8792 6554 8816 6556
rect 8872 6554 8896 6556
rect 8952 6554 8976 6556
rect 8712 6502 8722 6554
rect 8966 6502 8976 6554
rect 8712 6500 8736 6502
rect 8792 6500 8816 6502
rect 8872 6500 8896 6502
rect 8952 6500 8976 6502
rect 8656 6491 9032 6500
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9048 5658 9076 6258
rect 9140 5914 9168 11018
rect 9232 9110 9260 11018
rect 9310 10704 9366 10713
rect 9310 10639 9366 10648
rect 9324 9994 9352 10639
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9324 9518 9352 9930
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9220 9104 9272 9110
rect 9220 9046 9272 9052
rect 9324 8974 9352 9318
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9232 8634 9260 8910
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9416 8090 9444 12242
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9508 7970 9536 13126
rect 9416 7942 9536 7970
rect 9416 7868 9444 7942
rect 9232 7840 9444 7868
rect 9496 7880 9548 7886
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9232 5710 9260 7840
rect 9496 7822 9548 7828
rect 9404 6928 9456 6934
rect 9404 6870 9456 6876
rect 9220 5704 9272 5710
rect 9048 5630 9168 5658
rect 9220 5646 9272 5652
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 8656 5468 9032 5477
rect 8712 5466 8736 5468
rect 8792 5466 8816 5468
rect 8872 5466 8896 5468
rect 8952 5466 8976 5468
rect 8712 5414 8722 5466
rect 8966 5414 8976 5466
rect 8712 5412 8736 5414
rect 8792 5412 8816 5414
rect 8872 5412 8896 5414
rect 8952 5412 8976 5414
rect 8656 5403 9032 5412
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9048 4622 9076 5306
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 8656 4380 9032 4389
rect 8712 4378 8736 4380
rect 8792 4378 8816 4380
rect 8872 4378 8896 4380
rect 8952 4378 8976 4380
rect 8712 4326 8722 4378
rect 8966 4326 8976 4378
rect 8712 4324 8736 4326
rect 8792 4324 8816 4326
rect 8872 4324 8896 4326
rect 8952 4324 8976 4326
rect 8656 4315 9032 4324
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8588 3670 8616 3878
rect 9048 3738 9076 4218
rect 9140 3942 9168 5630
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9232 4078 9260 5510
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9324 3738 9352 5646
rect 9416 5234 9444 6870
rect 9508 6866 9536 7822
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9508 6322 9536 6802
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9404 4752 9456 4758
rect 9404 4694 9456 4700
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9416 3670 9444 4694
rect 9508 4570 9536 5510
rect 9600 4826 9628 14962
rect 9692 14618 9720 15846
rect 9784 15026 9812 16186
rect 9876 15502 9904 16390
rect 10520 15570 10548 16934
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10888 15502 10916 19110
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9876 14906 9904 15438
rect 9956 15428 10008 15434
rect 9956 15370 10008 15376
rect 9784 14878 9904 14906
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9784 14414 9812 14878
rect 9968 14822 9996 15370
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9680 13456 9732 13462
rect 9680 13398 9732 13404
rect 9692 11762 9720 13398
rect 9784 12714 9812 14350
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 9968 14006 9996 14282
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9770 12608 9826 12617
rect 9770 12543 9826 12552
rect 9784 11830 9812 12543
rect 9876 12238 9904 13942
rect 10796 13530 10824 14962
rect 10980 14822 11008 18702
rect 11072 15094 11100 19246
rect 11164 18850 11192 21286
rect 11256 21146 11284 21286
rect 11244 21140 11296 21146
rect 11244 21082 11296 21088
rect 11336 20868 11388 20874
rect 11336 20810 11388 20816
rect 11348 20602 11376 20810
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 11532 20398 11560 21508
rect 11612 21490 11664 21496
rect 11796 21480 11848 21486
rect 11796 21422 11848 21428
rect 11612 21344 11664 21350
rect 11612 21286 11664 21292
rect 11520 20392 11572 20398
rect 11520 20334 11572 20340
rect 11164 18822 11284 18850
rect 11532 18834 11560 20334
rect 11624 19854 11652 21286
rect 11808 20806 11836 21422
rect 11796 20800 11848 20806
rect 11796 20742 11848 20748
rect 11808 20534 11836 20742
rect 11796 20528 11848 20534
rect 11796 20470 11848 20476
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 11164 17882 11192 18702
rect 11256 18154 11284 18822
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11428 18624 11480 18630
rect 11428 18566 11480 18572
rect 11244 18148 11296 18154
rect 11244 18090 11296 18096
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11440 17202 11468 18566
rect 11612 17808 11664 17814
rect 11612 17750 11664 17756
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11520 17060 11572 17066
rect 11520 17002 11572 17008
rect 11532 16250 11560 17002
rect 11624 16794 11652 17750
rect 11716 17746 11744 19314
rect 11900 19310 11928 21626
rect 12084 19786 12112 21830
rect 12636 21554 12664 21966
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12452 21146 12480 21286
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12544 19854 12572 20878
rect 12636 20058 12664 21490
rect 13004 20058 13032 24142
rect 13916 23420 14292 23429
rect 13972 23418 13996 23420
rect 14052 23418 14076 23420
rect 14132 23418 14156 23420
rect 14212 23418 14236 23420
rect 13972 23366 13982 23418
rect 14226 23366 14236 23418
rect 13972 23364 13996 23366
rect 14052 23364 14076 23366
rect 14132 23364 14156 23366
rect 14212 23364 14236 23366
rect 13916 23355 14292 23364
rect 13916 22332 14292 22341
rect 13972 22330 13996 22332
rect 14052 22330 14076 22332
rect 14132 22330 14156 22332
rect 14212 22330 14236 22332
rect 13972 22278 13982 22330
rect 14226 22278 14236 22330
rect 13972 22276 13996 22278
rect 14052 22276 14076 22278
rect 14132 22276 14156 22278
rect 14212 22276 14236 22278
rect 13916 22267 14292 22276
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 13176 21956 13228 21962
rect 13176 21898 13228 21904
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12992 20052 13044 20058
rect 12992 19994 13044 20000
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12072 19780 12124 19786
rect 12072 19722 12124 19728
rect 13188 19378 13216 21898
rect 13268 21888 13320 21894
rect 13268 21830 13320 21836
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13280 19854 13308 21830
rect 13740 21622 13768 21830
rect 13728 21616 13780 21622
rect 13728 21558 13780 21564
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13740 20942 13768 21286
rect 13728 20936 13780 20942
rect 13728 20878 13780 20884
rect 13832 19854 13860 21830
rect 14292 21434 14320 21966
rect 14464 21888 14516 21894
rect 14464 21830 14516 21836
rect 14292 21406 14412 21434
rect 13916 21244 14292 21253
rect 13972 21242 13996 21244
rect 14052 21242 14076 21244
rect 14132 21242 14156 21244
rect 14212 21242 14236 21244
rect 13972 21190 13982 21242
rect 14226 21190 14236 21242
rect 13972 21188 13996 21190
rect 14052 21188 14076 21190
rect 14132 21188 14156 21190
rect 14212 21188 14236 21190
rect 13916 21179 14292 21188
rect 13916 20156 14292 20165
rect 13972 20154 13996 20156
rect 14052 20154 14076 20156
rect 14132 20154 14156 20156
rect 14212 20154 14236 20156
rect 13972 20102 13982 20154
rect 14226 20102 14236 20154
rect 13972 20100 13996 20102
rect 14052 20100 14076 20102
rect 14132 20100 14156 20102
rect 14212 20100 14236 20102
rect 13916 20091 14292 20100
rect 14384 20058 14412 21406
rect 14476 20602 14504 21830
rect 14568 21570 14596 24142
rect 14656 23964 15032 23973
rect 14712 23962 14736 23964
rect 14792 23962 14816 23964
rect 14872 23962 14896 23964
rect 14952 23962 14976 23964
rect 14712 23910 14722 23962
rect 14966 23910 14976 23962
rect 14712 23908 14736 23910
rect 14792 23908 14816 23910
rect 14872 23908 14896 23910
rect 14952 23908 14976 23910
rect 14656 23899 15032 23908
rect 14656 22876 15032 22885
rect 14712 22874 14736 22876
rect 14792 22874 14816 22876
rect 14872 22874 14896 22876
rect 14952 22874 14976 22876
rect 14712 22822 14722 22874
rect 14966 22822 14976 22874
rect 14712 22820 14736 22822
rect 14792 22820 14816 22822
rect 14872 22820 14896 22822
rect 14952 22820 14976 22822
rect 14656 22811 15032 22820
rect 15396 22094 15424 24142
rect 20656 23964 21032 23973
rect 20712 23962 20736 23964
rect 20792 23962 20816 23964
rect 20872 23962 20896 23964
rect 20952 23962 20976 23964
rect 20712 23910 20722 23962
rect 20966 23910 20976 23962
rect 20712 23908 20736 23910
rect 20792 23908 20816 23910
rect 20872 23908 20896 23910
rect 20952 23908 20976 23910
rect 20656 23899 21032 23908
rect 19916 23420 20292 23429
rect 19972 23418 19996 23420
rect 20052 23418 20076 23420
rect 20132 23418 20156 23420
rect 20212 23418 20236 23420
rect 19972 23366 19982 23418
rect 20226 23366 20236 23418
rect 19972 23364 19996 23366
rect 20052 23364 20076 23366
rect 20132 23364 20156 23366
rect 20212 23364 20236 23366
rect 19916 23355 20292 23364
rect 20656 22876 21032 22885
rect 20712 22874 20736 22876
rect 20792 22874 20816 22876
rect 20872 22874 20896 22876
rect 20952 22874 20976 22876
rect 20712 22822 20722 22874
rect 20966 22822 20976 22874
rect 20712 22820 20736 22822
rect 20792 22820 20816 22822
rect 20872 22820 20896 22822
rect 20952 22820 20976 22822
rect 20656 22811 21032 22820
rect 16488 22636 16540 22642
rect 16488 22578 16540 22584
rect 15396 22066 15700 22094
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 15476 21888 15528 21894
rect 15476 21830 15528 21836
rect 14656 21788 15032 21797
rect 14712 21786 14736 21788
rect 14792 21786 14816 21788
rect 14872 21786 14896 21788
rect 14952 21786 14976 21788
rect 14712 21734 14722 21786
rect 14966 21734 14976 21786
rect 14712 21732 14736 21734
rect 14792 21732 14816 21734
rect 14872 21732 14896 21734
rect 14952 21732 14976 21734
rect 14656 21723 15032 21732
rect 14568 21542 14688 21570
rect 14556 21480 14608 21486
rect 14556 21422 14608 21428
rect 14464 20596 14516 20602
rect 14464 20538 14516 20544
rect 14568 20346 14596 21422
rect 14660 20942 14688 21542
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 15200 21344 15252 21350
rect 15200 21286 15252 21292
rect 14752 21146 14780 21286
rect 14740 21140 14792 21146
rect 14740 21082 14792 21088
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14656 20700 15032 20709
rect 14712 20698 14736 20700
rect 14792 20698 14816 20700
rect 14872 20698 14896 20700
rect 14952 20698 14976 20700
rect 14712 20646 14722 20698
rect 14966 20646 14976 20698
rect 14712 20644 14736 20646
rect 14792 20644 14816 20646
rect 14872 20644 14896 20646
rect 14952 20644 14976 20646
rect 14656 20635 15032 20644
rect 15212 20466 15240 21286
rect 15304 21146 15332 21830
rect 15488 21554 15516 21830
rect 15476 21548 15528 21554
rect 15476 21490 15528 21496
rect 15384 21344 15436 21350
rect 15384 21286 15436 21292
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15396 20618 15424 21286
rect 15304 20590 15424 20618
rect 15304 20534 15332 20590
rect 15292 20528 15344 20534
rect 15292 20470 15344 20476
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 14476 20330 14596 20346
rect 14464 20324 14596 20330
rect 14516 20318 14596 20324
rect 14464 20266 14516 20272
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 14372 20052 14424 20058
rect 14372 19994 14424 20000
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 14384 19514 14412 19994
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 11888 19304 11940 19310
rect 11888 19246 11940 19252
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 11348 14822 11376 15982
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 10244 12102 10272 12378
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9692 8566 9720 9318
rect 9876 9178 9904 10066
rect 9864 9172 9916 9178
rect 9916 9132 9996 9160
rect 9864 9114 9916 9120
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9692 6730 9720 8502
rect 9876 7546 9904 8842
rect 9968 7818 9996 9132
rect 10244 8838 10272 12038
rect 11072 11898 11100 13874
rect 11164 13326 11192 14214
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 12646 11192 13126
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10336 9722 10364 10406
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10428 9586 10456 10406
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 9956 7812 10008 7818
rect 9956 7754 10008 7760
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9692 5370 9720 6666
rect 9876 6458 9904 7142
rect 9968 6730 9996 7142
rect 9956 6724 10008 6730
rect 9956 6666 10008 6672
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 9508 4542 9628 4570
rect 9600 4486 9628 4542
rect 9496 4480 9548 4486
rect 9496 4422 9548 4428
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 8576 3664 8628 3670
rect 8576 3606 8628 3612
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9508 3534 9536 4422
rect 9692 3534 9720 4966
rect 9784 4282 9812 5170
rect 9968 4690 9996 6258
rect 10060 5370 10088 8230
rect 10520 8022 10548 11698
rect 11256 11694 11284 13262
rect 11348 12986 11376 13806
rect 11624 13802 11652 14758
rect 11612 13796 11664 13802
rect 11612 13738 11664 13744
rect 11716 13682 11744 17138
rect 11808 15978 11836 18566
rect 11900 18222 11928 19246
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 11888 18216 11940 18222
rect 11888 18158 11940 18164
rect 11900 17678 11928 18158
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11900 16182 11928 17614
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 11796 15972 11848 15978
rect 11796 15914 11848 15920
rect 11900 14006 11928 16118
rect 11992 15706 12020 18566
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 12084 16250 12112 17546
rect 13188 17270 13216 18566
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 13280 17338 13308 18158
rect 13372 17882 13400 18702
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13176 17264 13228 17270
rect 13176 17206 13228 17212
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 12084 15162 12112 15438
rect 12348 15428 12400 15434
rect 12348 15370 12400 15376
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11992 14006 12020 14554
rect 12164 14340 12216 14346
rect 12164 14282 12216 14288
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 11440 13654 11744 13682
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11348 12646 11376 12786
rect 11440 12714 11468 13654
rect 11610 13424 11666 13433
rect 11610 13359 11666 13368
rect 11624 13326 11652 13359
rect 11900 13326 11928 13942
rect 12176 13938 12204 14282
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11428 12708 11480 12714
rect 11428 12650 11480 12656
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10612 9586 10640 10134
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10508 8016 10560 8022
rect 10508 7958 10560 7964
rect 10704 7954 10732 9862
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10796 7886 10824 11086
rect 11164 11082 11192 11494
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11164 10130 11192 11018
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11242 9616 11298 9625
rect 11242 9551 11298 9560
rect 11256 9382 11284 9551
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10324 7744 10376 7750
rect 11348 7698 11376 12038
rect 10324 7686 10376 7692
rect 10336 6458 10364 7686
rect 11256 7670 11376 7698
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9876 4146 9904 4626
rect 10060 4554 10088 5306
rect 10244 5030 10272 6258
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10336 4554 10364 5850
rect 10416 5636 10468 5642
rect 10416 5578 10468 5584
rect 10428 5302 10456 5578
rect 10520 5302 10548 6938
rect 11256 6769 11284 7670
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 11242 6760 11298 6769
rect 11242 6695 11298 6704
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11072 5710 11100 6598
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 10416 5296 10468 5302
rect 10416 5238 10468 5244
rect 10508 5296 10560 5302
rect 10508 5238 10560 5244
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10048 4548 10100 4554
rect 10048 4490 10100 4496
rect 10324 4548 10376 4554
rect 10324 4490 10376 4496
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 10704 4078 10732 4966
rect 10796 4146 10824 5646
rect 11256 4146 11284 6598
rect 11348 6458 11376 7482
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11348 5710 11376 6054
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 11072 3534 11100 3946
rect 11348 3738 11376 5102
rect 11440 4622 11468 12650
rect 11532 10538 11560 12786
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11624 11762 11652 12718
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11716 11354 11744 11698
rect 11808 11558 11836 12582
rect 12360 12374 12388 15370
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 12900 14000 12952 14006
rect 12900 13942 12952 13948
rect 12912 13530 12940 13942
rect 13004 13530 13032 14010
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 13188 13394 13216 16390
rect 13280 16250 13308 17274
rect 13556 16522 13584 18566
rect 13740 17678 13768 19450
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 13916 19068 14292 19077
rect 13972 19066 13996 19068
rect 14052 19066 14076 19068
rect 14132 19066 14156 19068
rect 14212 19066 14236 19068
rect 13972 19014 13982 19066
rect 14226 19014 14236 19066
rect 13972 19012 13996 19014
rect 14052 19012 14076 19014
rect 14132 19012 14156 19014
rect 14212 19012 14236 19014
rect 13916 19003 14292 19012
rect 13820 18692 13872 18698
rect 13820 18634 13872 18640
rect 14004 18692 14056 18698
rect 14004 18634 14056 18640
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13648 17338 13676 17478
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 13832 16454 13860 18634
rect 14016 18426 14044 18634
rect 14280 18624 14332 18630
rect 14280 18566 14332 18572
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 14292 18170 14320 18566
rect 14384 18426 14412 19314
rect 14476 18766 14504 19790
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14568 19394 14596 19654
rect 14656 19612 15032 19621
rect 14712 19610 14736 19612
rect 14792 19610 14816 19612
rect 14872 19610 14896 19612
rect 14952 19610 14976 19612
rect 14712 19558 14722 19610
rect 14966 19558 14976 19610
rect 14712 19556 14736 19558
rect 14792 19556 14816 19558
rect 14872 19556 14896 19558
rect 14952 19556 14976 19558
rect 14656 19547 15032 19556
rect 14922 19408 14978 19417
rect 14568 19366 14688 19394
rect 14556 19304 14608 19310
rect 14556 19246 14608 19252
rect 14568 18970 14596 19246
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14660 18834 14688 19366
rect 15120 19378 15148 20198
rect 15292 19984 15344 19990
rect 15292 19926 15344 19932
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15212 19514 15240 19790
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 14922 19343 14978 19352
rect 15108 19372 15160 19378
rect 14936 19174 14964 19343
rect 15108 19314 15160 19320
rect 14924 19168 14976 19174
rect 14924 19110 14976 19116
rect 14648 18828 14700 18834
rect 14648 18770 14700 18776
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14292 18142 14412 18170
rect 13916 17980 14292 17989
rect 13972 17978 13996 17980
rect 14052 17978 14076 17980
rect 14132 17978 14156 17980
rect 14212 17978 14236 17980
rect 13972 17926 13982 17978
rect 14226 17926 14236 17978
rect 13972 17924 13996 17926
rect 14052 17924 14076 17926
rect 14132 17924 14156 17926
rect 14212 17924 14236 17926
rect 13916 17915 14292 17924
rect 14384 17678 14412 18142
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14384 17270 14412 17478
rect 14372 17264 14424 17270
rect 14372 17206 14424 17212
rect 13916 16892 14292 16901
rect 13972 16890 13996 16892
rect 14052 16890 14076 16892
rect 14132 16890 14156 16892
rect 14212 16890 14236 16892
rect 13972 16838 13982 16890
rect 14226 16838 14236 16890
rect 13972 16836 13996 16838
rect 14052 16836 14076 16838
rect 14132 16836 14156 16838
rect 14212 16836 14236 16838
rect 13916 16827 14292 16836
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13832 16114 13860 16390
rect 14384 16250 14412 16594
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 13912 16176 13964 16182
rect 13912 16118 13964 16124
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13728 16040 13780 16046
rect 13924 15994 13952 16118
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 13728 15982 13780 15988
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 13464 15094 13492 15846
rect 13740 15706 13768 15982
rect 13832 15966 13952 15994
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13832 15586 13860 15966
rect 13916 15804 14292 15813
rect 13972 15802 13996 15804
rect 14052 15802 14076 15804
rect 14132 15802 14156 15804
rect 14212 15802 14236 15804
rect 13972 15750 13982 15802
rect 14226 15750 14236 15802
rect 13972 15748 13996 15750
rect 14052 15748 14076 15750
rect 14132 15748 14156 15750
rect 14212 15748 14236 15750
rect 13916 15739 14292 15748
rect 13832 15558 13952 15586
rect 14384 15570 14412 16050
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13452 15088 13504 15094
rect 13452 15030 13504 15036
rect 13832 15026 13860 15302
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13924 14906 13952 15558
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 14372 15156 14424 15162
rect 14372 15098 14424 15104
rect 13832 14878 13952 14906
rect 13832 14550 13860 14878
rect 14384 14822 14412 15098
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 13916 14716 14292 14725
rect 13972 14714 13996 14716
rect 14052 14714 14076 14716
rect 14132 14714 14156 14716
rect 14212 14714 14236 14716
rect 13972 14662 13982 14714
rect 14226 14662 14236 14714
rect 13972 14660 13996 14662
rect 14052 14660 14076 14662
rect 14132 14660 14156 14662
rect 14212 14660 14236 14662
rect 13916 14651 14292 14660
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13372 14074 13400 14350
rect 14188 14340 14240 14346
rect 14188 14282 14240 14288
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12348 12368 12400 12374
rect 12348 12310 12400 12316
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11624 10674 11652 11222
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11520 10532 11572 10538
rect 11520 10474 11572 10480
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11532 9586 11560 9998
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11532 7478 11560 9522
rect 11520 7472 11572 7478
rect 11520 7414 11572 7420
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11336 3732 11388 3738
rect 11336 3674 11388 3680
rect 11532 3670 11560 7278
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11624 3534 11652 9862
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11716 6254 11744 9454
rect 11808 7546 11836 9998
rect 11900 9625 11928 12106
rect 12820 11830 12848 12922
rect 13372 12238 13400 14010
rect 13556 14006 13584 14214
rect 14200 14074 14228 14282
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 13820 13932 13872 13938
rect 13740 13892 13820 13920
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13464 12442 13492 13262
rect 13636 12844 13688 12850
rect 13556 12804 13636 12832
rect 13556 12442 13584 12804
rect 13636 12786 13688 12792
rect 13740 12730 13768 13892
rect 13820 13874 13872 13880
rect 13820 13796 13872 13802
rect 13820 13738 13872 13744
rect 13832 13512 13860 13738
rect 13916 13628 14292 13637
rect 13972 13626 13996 13628
rect 14052 13626 14076 13628
rect 14132 13626 14156 13628
rect 14212 13626 14236 13628
rect 13972 13574 13982 13626
rect 14226 13574 14236 13626
rect 13972 13572 13996 13574
rect 14052 13572 14076 13574
rect 14132 13572 14156 13574
rect 14212 13572 14236 13574
rect 13916 13563 14292 13572
rect 14384 13530 14412 14758
rect 14372 13524 14424 13530
rect 13832 13484 13952 13512
rect 13820 13252 13872 13258
rect 13820 13194 13872 13200
rect 13648 12702 13768 12730
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13648 12322 13676 12702
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13464 12306 13676 12322
rect 13452 12300 13676 12306
rect 13504 12294 13676 12300
rect 13452 12242 13504 12248
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12544 10062 12572 10406
rect 12820 10062 12848 11290
rect 13004 11150 13032 11494
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13280 11150 13308 11290
rect 13648 11150 13676 12038
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13740 10674 13768 12582
rect 13832 10810 13860 13194
rect 13924 12850 13952 13484
rect 14372 13466 14424 13472
rect 14370 13424 14426 13433
rect 14370 13359 14426 13368
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 14278 12744 14334 12753
rect 14278 12679 14280 12688
rect 14332 12679 14334 12688
rect 14280 12650 14332 12656
rect 14384 12646 14412 13359
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 13916 12540 14292 12549
rect 13972 12538 13996 12540
rect 14052 12538 14076 12540
rect 14132 12538 14156 12540
rect 14212 12538 14236 12540
rect 13972 12486 13982 12538
rect 14226 12486 14236 12538
rect 13972 12484 13996 12486
rect 14052 12484 14076 12486
rect 14132 12484 14156 12486
rect 14212 12484 14236 12486
rect 13916 12475 14292 12484
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 13916 11452 14292 11461
rect 13972 11450 13996 11452
rect 14052 11450 14076 11452
rect 14132 11450 14156 11452
rect 14212 11450 14236 11452
rect 13972 11398 13982 11450
rect 14226 11398 14236 11450
rect 13972 11396 13996 11398
rect 14052 11396 14076 11398
rect 14132 11396 14156 11398
rect 14212 11396 14236 11398
rect 13916 11387 14292 11396
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13648 10266 13676 10610
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 12532 10056 12584 10062
rect 12808 10056 12860 10062
rect 12532 9998 12584 10004
rect 12622 10024 12678 10033
rect 12808 9998 12860 10004
rect 12622 9959 12624 9968
rect 12676 9959 12678 9968
rect 12624 9930 12676 9936
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 11980 9648 12032 9654
rect 11886 9616 11942 9625
rect 11980 9590 12032 9596
rect 12544 9602 12572 9862
rect 11886 9551 11942 9560
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11716 5098 11744 5510
rect 11704 5092 11756 5098
rect 11704 5034 11756 5040
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 8656 3292 9032 3301
rect 8712 3290 8736 3292
rect 8792 3290 8816 3292
rect 8872 3290 8896 3292
rect 8952 3290 8976 3292
rect 8712 3238 8722 3290
rect 8966 3238 8976 3290
rect 8712 3236 8736 3238
rect 8792 3236 8816 3238
rect 8872 3236 8896 3238
rect 8952 3236 8976 3238
rect 8656 3227 9032 3236
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 7916 2748 8292 2757
rect 7972 2746 7996 2748
rect 8052 2746 8076 2748
rect 8132 2746 8156 2748
rect 8212 2746 8236 2748
rect 7972 2694 7982 2746
rect 8226 2694 8236 2746
rect 7972 2692 7996 2694
rect 8052 2692 8076 2694
rect 8132 2692 8156 2694
rect 8212 2692 8236 2694
rect 7916 2683 8292 2692
rect 6276 2576 6328 2582
rect 6276 2518 6328 2524
rect 7116 2514 7236 2530
rect 7116 2508 7248 2514
rect 7116 2502 7196 2508
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 2656 2204 3032 2213
rect 2712 2202 2736 2204
rect 2792 2202 2816 2204
rect 2872 2202 2896 2204
rect 2952 2202 2976 2204
rect 2712 2150 2722 2202
rect 2966 2150 2976 2202
rect 2712 2148 2736 2150
rect 2792 2148 2816 2150
rect 2872 2148 2896 2150
rect 2952 2148 2976 2150
rect 2656 2139 3032 2148
rect 7116 800 7144 2502
rect 7196 2450 7248 2456
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 7760 800 7788 2314
rect 8656 2204 9032 2213
rect 8712 2202 8736 2204
rect 8792 2202 8816 2204
rect 8872 2202 8896 2204
rect 8952 2202 8976 2204
rect 8712 2150 8722 2202
rect 8966 2150 8976 2202
rect 8712 2148 8736 2150
rect 8792 2148 8816 2150
rect 8872 2148 8896 2150
rect 8952 2148 8976 2150
rect 8656 2139 9032 2148
rect 10428 1306 10456 2382
rect 10336 1278 10456 1306
rect 10336 800 10364 1278
rect 10980 800 11008 2926
rect 11808 2514 11836 7278
rect 11900 7274 11928 9318
rect 11992 9178 12020 9590
rect 12544 9574 12664 9602
rect 12532 9512 12584 9518
rect 12438 9480 12494 9489
rect 12532 9454 12584 9460
rect 12438 9415 12494 9424
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11992 8022 12020 9114
rect 12452 8498 12480 9415
rect 12544 9178 12572 9454
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 12162 7984 12218 7993
rect 11888 7268 11940 7274
rect 11888 7210 11940 7216
rect 11992 4162 12020 7958
rect 12162 7919 12218 7928
rect 12176 7886 12204 7919
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 12084 7410 12112 7686
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 11900 4146 12020 4162
rect 11888 4140 12020 4146
rect 11940 4134 12020 4140
rect 11888 4082 11940 4088
rect 11992 3534 12020 4134
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 12268 2446 12296 4422
rect 12452 3738 12480 6734
rect 12636 6338 12664 9574
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 12992 9444 13044 9450
rect 12992 9386 13044 9392
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12820 9178 12848 9318
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12728 7410 12756 7754
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12544 6310 12664 6338
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12544 2446 12572 6310
rect 12728 5914 12756 7346
rect 13004 5914 13032 9386
rect 13464 7342 13492 9522
rect 13832 8974 13860 10610
rect 14108 10606 14136 11154
rect 14280 11076 14332 11082
rect 14280 11018 14332 11024
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14292 10554 14320 11018
rect 14384 10674 14412 12038
rect 14476 11665 14504 18226
rect 14568 16114 14596 18702
rect 14656 18524 15032 18533
rect 14712 18522 14736 18524
rect 14792 18522 14816 18524
rect 14872 18522 14896 18524
rect 14952 18522 14976 18524
rect 14712 18470 14722 18522
rect 14966 18470 14976 18522
rect 14712 18468 14736 18470
rect 14792 18468 14816 18470
rect 14872 18468 14896 18470
rect 14952 18468 14976 18470
rect 14656 18459 15032 18468
rect 15108 18420 15160 18426
rect 15108 18362 15160 18368
rect 14648 18148 14700 18154
rect 14648 18090 14700 18096
rect 14660 17882 14688 18090
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 14752 17542 14780 18022
rect 15120 17610 15148 18362
rect 15212 18154 15240 18770
rect 15200 18148 15252 18154
rect 15200 18090 15252 18096
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14656 17436 15032 17445
rect 14712 17434 14736 17436
rect 14792 17434 14816 17436
rect 14872 17434 14896 17436
rect 14952 17434 14976 17436
rect 14712 17382 14722 17434
rect 14966 17382 14976 17434
rect 14712 17380 14736 17382
rect 14792 17380 14816 17382
rect 14872 17380 14896 17382
rect 14952 17380 14976 17382
rect 14656 17371 15032 17380
rect 15304 17202 15332 19926
rect 15488 19854 15516 21490
rect 15568 21480 15620 21486
rect 15568 21422 15620 21428
rect 15580 21146 15608 21422
rect 15568 21140 15620 21146
rect 15568 21082 15620 21088
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 15488 18902 15516 19790
rect 15580 19417 15608 20742
rect 15566 19408 15622 19417
rect 15566 19343 15622 19352
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15672 17338 15700 22066
rect 16304 21344 16356 21350
rect 16304 21286 16356 21292
rect 16316 20942 16344 21286
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 16500 20262 16528 22578
rect 19916 22332 20292 22341
rect 19972 22330 19996 22332
rect 20052 22330 20076 22332
rect 20132 22330 20156 22332
rect 20212 22330 20236 22332
rect 19972 22278 19982 22330
rect 20226 22278 20236 22330
rect 19972 22276 19996 22278
rect 20052 22276 20076 22278
rect 20132 22276 20156 22278
rect 20212 22276 20236 22278
rect 19916 22267 20292 22276
rect 20656 21788 21032 21797
rect 20712 21786 20736 21788
rect 20792 21786 20816 21788
rect 20872 21786 20896 21788
rect 20952 21786 20976 21788
rect 20712 21734 20722 21786
rect 20966 21734 20976 21786
rect 20712 21732 20736 21734
rect 20792 21732 20816 21734
rect 20872 21732 20896 21734
rect 20952 21732 20976 21734
rect 20656 21723 21032 21732
rect 17224 21480 17276 21486
rect 17224 21422 17276 21428
rect 18144 21480 18196 21486
rect 18144 21422 18196 21428
rect 16672 21344 16724 21350
rect 16672 21286 16724 21292
rect 16684 20398 16712 21286
rect 17236 20602 17264 21422
rect 17776 20936 17828 20942
rect 17776 20878 17828 20884
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 16672 20392 16724 20398
rect 16672 20334 16724 20340
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17408 20392 17460 20398
rect 17408 20334 17460 20340
rect 16488 20256 16540 20262
rect 16488 20198 16540 20204
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16684 19242 16712 20198
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 16764 19440 16816 19446
rect 16764 19382 16816 19388
rect 16672 19236 16724 19242
rect 16672 19178 16724 19184
rect 16776 18290 16804 19382
rect 16856 18352 16908 18358
rect 16856 18294 16908 18300
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 14656 16348 15032 16357
rect 14712 16346 14736 16348
rect 14792 16346 14816 16348
rect 14872 16346 14896 16348
rect 14952 16346 14976 16348
rect 14712 16294 14722 16346
rect 14966 16294 14976 16346
rect 14712 16292 14736 16294
rect 14792 16292 14816 16294
rect 14872 16292 14896 16294
rect 14952 16292 14976 16294
rect 14656 16283 15032 16292
rect 15856 16250 15884 16526
rect 15936 16516 15988 16522
rect 15936 16458 15988 16464
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14568 12442 14596 15302
rect 14656 15260 15032 15269
rect 14712 15258 14736 15260
rect 14792 15258 14816 15260
rect 14872 15258 14896 15260
rect 14952 15258 14976 15260
rect 14712 15206 14722 15258
rect 14966 15206 14976 15258
rect 14712 15204 14736 15206
rect 14792 15204 14816 15206
rect 14872 15204 14896 15206
rect 14952 15204 14976 15206
rect 14656 15195 15032 15204
rect 14656 14172 15032 14181
rect 14712 14170 14736 14172
rect 14792 14170 14816 14172
rect 14872 14170 14896 14172
rect 14952 14170 14976 14172
rect 14712 14118 14722 14170
rect 14966 14118 14976 14170
rect 14712 14116 14736 14118
rect 14792 14116 14816 14118
rect 14872 14116 14896 14118
rect 14952 14116 14976 14118
rect 14656 14107 15032 14116
rect 15120 14006 15148 15846
rect 15200 15428 15252 15434
rect 15200 15370 15252 15376
rect 15212 14482 15240 15370
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15108 14000 15160 14006
rect 15108 13942 15160 13948
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14844 13394 14872 13670
rect 14832 13388 14884 13394
rect 14832 13330 14884 13336
rect 15304 13274 15332 16050
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15396 14414 15424 15642
rect 15488 15434 15516 15642
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 15120 13246 15332 13274
rect 14656 13084 15032 13093
rect 14712 13082 14736 13084
rect 14792 13082 14816 13084
rect 14872 13082 14896 13084
rect 14952 13082 14976 13084
rect 14712 13030 14722 13082
rect 14966 13030 14976 13082
rect 14712 13028 14736 13030
rect 14792 13028 14816 13030
rect 14872 13028 14896 13030
rect 14952 13028 14976 13030
rect 14656 13019 15032 13028
rect 15120 12850 15148 13246
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 14556 12436 14608 12442
rect 14556 12378 14608 12384
rect 14656 11996 15032 12005
rect 14712 11994 14736 11996
rect 14792 11994 14816 11996
rect 14872 11994 14896 11996
rect 14952 11994 14976 11996
rect 14712 11942 14722 11994
rect 14966 11942 14976 11994
rect 14712 11940 14736 11942
rect 14792 11940 14816 11942
rect 14872 11940 14896 11942
rect 14952 11940 14976 11942
rect 14656 11931 15032 11940
rect 15108 11824 15160 11830
rect 15108 11766 15160 11772
rect 14462 11656 14518 11665
rect 14462 11591 14518 11600
rect 15120 11150 15148 11766
rect 15212 11370 15240 12854
rect 15304 12442 15332 13126
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15212 11342 15332 11370
rect 15304 11286 15332 11342
rect 15292 11280 15344 11286
rect 15292 11222 15344 11228
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 14656 10908 15032 10917
rect 14712 10906 14736 10908
rect 14792 10906 14816 10908
rect 14872 10906 14896 10908
rect 14952 10906 14976 10908
rect 14712 10854 14722 10906
rect 14966 10854 14976 10906
rect 14712 10852 14736 10854
rect 14792 10852 14816 10854
rect 14872 10852 14896 10854
rect 14952 10852 14976 10854
rect 14656 10843 15032 10852
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14292 10526 14412 10554
rect 13916 10364 14292 10373
rect 13972 10362 13996 10364
rect 14052 10362 14076 10364
rect 14132 10362 14156 10364
rect 14212 10362 14236 10364
rect 13972 10310 13982 10362
rect 14226 10310 14236 10362
rect 13972 10308 13996 10310
rect 14052 10308 14076 10310
rect 14132 10308 14156 10310
rect 14212 10308 14236 10310
rect 13916 10299 14292 10308
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 14108 9586 14136 9930
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14200 9382 14228 10066
rect 14384 9874 14412 10526
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14292 9846 14412 9874
rect 14292 9654 14320 9846
rect 14476 9722 14504 10406
rect 14660 10010 14688 10610
rect 14568 9982 14688 10010
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 13916 9276 14292 9285
rect 13972 9274 13996 9276
rect 14052 9274 14076 9276
rect 14132 9274 14156 9276
rect 14212 9274 14236 9276
rect 13972 9222 13982 9274
rect 14226 9222 14236 9274
rect 13972 9220 13996 9222
rect 14052 9220 14076 9222
rect 14132 9220 14156 9222
rect 14212 9220 14236 9222
rect 13916 9211 14292 9220
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 13556 7546 13584 8842
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12636 5302 12664 5782
rect 12624 5296 12676 5302
rect 12624 5238 12676 5244
rect 12636 4214 12664 5238
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 12912 3942 12940 5170
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 13004 4622 13032 4966
rect 13096 4826 13124 7142
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 13188 4214 13216 4558
rect 13176 4208 13228 4214
rect 13176 4150 13228 4156
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 13372 2446 13400 6598
rect 13556 5370 13584 7142
rect 13648 6458 13676 7754
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 13556 4622 13584 5306
rect 13648 5250 13676 6258
rect 13740 5846 13768 8366
rect 13832 6798 13860 8774
rect 13924 8634 13952 8910
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 14200 8566 14228 8910
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 13916 8188 14292 8197
rect 13972 8186 13996 8188
rect 14052 8186 14076 8188
rect 14132 8186 14156 8188
rect 14212 8186 14236 8188
rect 13972 8134 13982 8186
rect 14226 8134 14236 8186
rect 13972 8132 13996 8134
rect 14052 8132 14076 8134
rect 14132 8132 14156 8134
rect 14212 8132 14236 8134
rect 13916 8123 14292 8132
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14200 7290 14228 7686
rect 14292 7546 14320 8026
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14384 7410 14412 9658
rect 14568 9058 14596 9982
rect 14656 9820 15032 9829
rect 14712 9818 14736 9820
rect 14792 9818 14816 9820
rect 14872 9818 14896 9820
rect 14952 9818 14976 9820
rect 14712 9766 14722 9818
rect 14966 9766 14976 9818
rect 14712 9764 14736 9766
rect 14792 9764 14816 9766
rect 14872 9764 14896 9766
rect 14952 9764 14976 9766
rect 14656 9755 15032 9764
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 14476 9030 14596 9058
rect 14476 8090 14504 9030
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14200 7262 14412 7290
rect 13916 7100 14292 7109
rect 13972 7098 13996 7100
rect 14052 7098 14076 7100
rect 14132 7098 14156 7100
rect 14212 7098 14236 7100
rect 13972 7046 13982 7098
rect 14226 7046 14236 7098
rect 13972 7044 13996 7046
rect 14052 7044 14076 7046
rect 14132 7044 14156 7046
rect 14212 7044 14236 7046
rect 13916 7035 14292 7044
rect 14384 6798 14412 7262
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 13832 5370 13860 6258
rect 14108 6254 14136 6734
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 13916 6012 14292 6021
rect 13972 6010 13996 6012
rect 14052 6010 14076 6012
rect 14132 6010 14156 6012
rect 14212 6010 14236 6012
rect 13972 5958 13982 6010
rect 14226 5958 14236 6010
rect 13972 5956 13996 5958
rect 14052 5956 14076 5958
rect 14132 5956 14156 5958
rect 14212 5956 14236 5958
rect 13916 5947 14292 5956
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14200 5370 14228 5646
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 13648 5222 13860 5250
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13556 3534 13584 4558
rect 13740 4282 13768 5102
rect 13832 4826 13860 5222
rect 13916 4924 14292 4933
rect 13972 4922 13996 4924
rect 14052 4922 14076 4924
rect 14132 4922 14156 4924
rect 14212 4922 14236 4924
rect 13972 4870 13982 4922
rect 14226 4870 14236 4922
rect 13972 4868 13996 4870
rect 14052 4868 14076 4870
rect 14132 4868 14156 4870
rect 14212 4868 14236 4870
rect 13916 4859 14292 4868
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 14384 4010 14412 6054
rect 14476 5166 14504 7686
rect 14568 5234 14596 8842
rect 14660 8838 14688 9590
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14656 8732 15032 8741
rect 14712 8730 14736 8732
rect 14792 8730 14816 8732
rect 14872 8730 14896 8732
rect 14952 8730 14976 8732
rect 14712 8678 14722 8730
rect 14966 8678 14976 8730
rect 14712 8676 14736 8678
rect 14792 8676 14816 8678
rect 14872 8676 14896 8678
rect 14952 8676 14976 8678
rect 14656 8667 15032 8676
rect 15120 8514 15148 11086
rect 15304 8634 15332 11222
rect 15396 11082 15424 13398
rect 15476 13252 15528 13258
rect 15476 13194 15528 13200
rect 15488 11354 15516 13194
rect 15764 11898 15792 14758
rect 15948 13530 15976 16458
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16132 15706 16160 15846
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 15948 12434 15976 13466
rect 16224 12714 16252 16390
rect 16500 15570 16528 17478
rect 16868 17338 16896 18294
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16960 17882 16988 18226
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 17052 17338 17080 19722
rect 17236 19378 17264 20334
rect 17420 19446 17448 20334
rect 17788 20058 17816 20878
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 18064 20466 18092 20742
rect 18156 20534 18184 21422
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 18420 20936 18472 20942
rect 18420 20878 18472 20884
rect 18144 20528 18196 20534
rect 18144 20470 18196 20476
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 17776 20052 17828 20058
rect 17776 19994 17828 20000
rect 18052 19780 18104 19786
rect 18052 19722 18104 19728
rect 17408 19440 17460 19446
rect 17408 19382 17460 19388
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17972 17814 18000 18566
rect 18064 18426 18092 19722
rect 18156 19718 18184 20470
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 18432 19378 18460 20878
rect 18800 20534 18828 21286
rect 19916 21244 20292 21253
rect 19972 21242 19996 21244
rect 20052 21242 20076 21244
rect 20132 21242 20156 21244
rect 20212 21242 20236 21244
rect 19972 21190 19982 21242
rect 20226 21190 20236 21242
rect 19972 21188 19996 21190
rect 20052 21188 20076 21190
rect 20132 21188 20156 21190
rect 20212 21188 20236 21190
rect 19916 21179 20292 21188
rect 19524 20868 19576 20874
rect 19524 20810 19576 20816
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 18788 20528 18840 20534
rect 18788 20470 18840 20476
rect 19352 19854 19380 20742
rect 19536 19854 19564 20810
rect 20656 20700 21032 20709
rect 20712 20698 20736 20700
rect 20792 20698 20816 20700
rect 20872 20698 20896 20700
rect 20952 20698 20976 20700
rect 20712 20646 20722 20698
rect 20966 20646 20976 20698
rect 20712 20644 20736 20646
rect 20792 20644 20816 20646
rect 20872 20644 20896 20646
rect 20952 20644 20976 20646
rect 20656 20635 21032 20644
rect 19800 20256 19852 20262
rect 19800 20198 19852 20204
rect 21456 20256 21508 20262
rect 21456 20198 21508 20204
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 18144 19372 18196 19378
rect 18144 19314 18196 19320
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 18156 18426 18184 19314
rect 18236 19304 18288 19310
rect 18236 19246 18288 19252
rect 18248 18970 18276 19246
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 18052 18420 18104 18426
rect 18052 18362 18104 18368
rect 18144 18420 18196 18426
rect 18144 18362 18196 18368
rect 18524 17882 18552 19790
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18972 19712 19024 19718
rect 18972 19654 19024 19660
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 18708 18834 18736 19654
rect 18984 18834 19012 19654
rect 19352 19378 19380 19654
rect 19524 19440 19576 19446
rect 19524 19382 19576 19388
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 18696 18828 18748 18834
rect 18696 18770 18748 18776
rect 18972 18828 19024 18834
rect 18972 18770 19024 18776
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18892 17814 18920 18702
rect 17960 17808 18012 17814
rect 17960 17750 18012 17756
rect 18880 17808 18932 17814
rect 18880 17750 18932 17756
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16580 15904 16632 15910
rect 16580 15846 16632 15852
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16592 15026 16620 15846
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 16316 14618 16344 14894
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16304 14612 16356 14618
rect 16304 14554 16356 14560
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16408 14074 16436 14214
rect 16500 14074 16528 14758
rect 16684 14226 16712 16050
rect 16684 14198 16804 14226
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16396 13456 16448 13462
rect 16396 13398 16448 13404
rect 16212 12708 16264 12714
rect 16212 12650 16264 12656
rect 16408 12434 16436 13398
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 15948 12406 16068 12434
rect 16040 12238 16068 12406
rect 16316 12406 16436 12434
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15580 10810 15608 11698
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 16132 10674 16160 12038
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 15568 10056 15620 10062
rect 15474 10024 15530 10033
rect 15568 9998 15620 10004
rect 15474 9959 15530 9968
rect 15488 9654 15516 9959
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 14936 8486 15148 8514
rect 15396 8498 15424 9318
rect 15384 8492 15436 8498
rect 14936 8242 14964 8486
rect 15384 8434 15436 8440
rect 15016 8424 15068 8430
rect 15068 8372 15240 8378
rect 15016 8366 15240 8372
rect 15028 8350 15240 8366
rect 14936 8214 15148 8242
rect 14656 7644 15032 7653
rect 14712 7642 14736 7644
rect 14792 7642 14816 7644
rect 14872 7642 14896 7644
rect 14952 7642 14976 7644
rect 14712 7590 14722 7642
rect 14966 7590 14976 7642
rect 14712 7588 14736 7590
rect 14792 7588 14816 7590
rect 14872 7588 14896 7590
rect 14952 7588 14976 7590
rect 14656 7579 15032 7588
rect 14656 6556 15032 6565
rect 14712 6554 14736 6556
rect 14792 6554 14816 6556
rect 14872 6554 14896 6556
rect 14952 6554 14976 6556
rect 14712 6502 14722 6554
rect 14966 6502 14976 6554
rect 14712 6500 14736 6502
rect 14792 6500 14816 6502
rect 14872 6500 14896 6502
rect 14952 6500 14976 6502
rect 14656 6491 15032 6500
rect 15120 5642 15148 8214
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 14656 5468 15032 5477
rect 14712 5466 14736 5468
rect 14792 5466 14816 5468
rect 14872 5466 14896 5468
rect 14952 5466 14976 5468
rect 14712 5414 14722 5466
rect 14966 5414 14976 5466
rect 14712 5412 14736 5414
rect 14792 5412 14816 5414
rect 14872 5412 14896 5414
rect 14952 5412 14976 5414
rect 14656 5403 15032 5412
rect 15212 5234 15240 8350
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15304 5370 15332 6394
rect 15396 5574 15424 8434
rect 15580 7546 15608 9998
rect 16224 8634 16252 11494
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15764 6662 15792 8434
rect 16132 8362 16160 8570
rect 16316 8498 16344 12406
rect 16684 12170 16712 12718
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16776 11558 16804 14198
rect 16868 12986 16896 17138
rect 17040 16244 17092 16250
rect 16960 16204 17040 16232
rect 16960 15570 16988 16204
rect 17040 16186 17092 16192
rect 17880 16182 17908 17274
rect 18064 16658 18092 17614
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 18156 17338 18184 17478
rect 18144 17332 18196 17338
rect 18144 17274 18196 17280
rect 18512 16992 18564 16998
rect 18512 16934 18564 16940
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 18052 16652 18104 16658
rect 18052 16594 18104 16600
rect 17868 16176 17920 16182
rect 17868 16118 17920 16124
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 17040 15632 17092 15638
rect 17040 15574 17092 15580
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16960 12850 16988 15506
rect 17052 14618 17080 15574
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 17052 13938 17080 14554
rect 17144 14414 17172 15642
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 17604 15094 17632 15438
rect 17592 15088 17644 15094
rect 17592 15030 17644 15036
rect 17972 15026 18000 15846
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17684 15020 17736 15026
rect 17684 14962 17736 14968
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17236 14074 17264 14962
rect 17696 14074 17724 14962
rect 18064 14906 18092 16594
rect 18432 16590 18460 16730
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 18236 16448 18288 16454
rect 18236 16390 18288 16396
rect 18144 15428 18196 15434
rect 18144 15370 18196 15376
rect 17972 14878 18092 14906
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17684 14068 17736 14074
rect 17684 14010 17736 14016
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17132 13796 17184 13802
rect 17132 13738 17184 13744
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17052 12986 17080 13262
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 17144 12730 17172 13738
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 16868 12714 17172 12730
rect 16856 12708 17172 12714
rect 16908 12702 17172 12708
rect 16856 12650 16908 12656
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 16684 10826 16712 11154
rect 16592 10810 16712 10826
rect 16580 10804 16712 10810
rect 16632 10798 16712 10804
rect 16580 10746 16632 10752
rect 16672 10736 16724 10742
rect 16672 10678 16724 10684
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16592 9674 16620 10542
rect 16408 9654 16620 9674
rect 16684 9654 16712 10678
rect 16396 9648 16620 9654
rect 16448 9646 16620 9648
rect 16672 9648 16724 9654
rect 16396 9590 16448 9596
rect 16672 9590 16724 9596
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16408 8090 16436 8230
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15488 5642 15516 6054
rect 15672 5914 15700 6054
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15476 5636 15528 5642
rect 15476 5578 15528 5584
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15672 5370 15700 5646
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14568 4622 14596 5170
rect 15856 5166 15884 7346
rect 15948 6458 15976 7822
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 16040 5370 16068 7822
rect 16304 7812 16356 7818
rect 16304 7754 16356 7760
rect 16120 7744 16172 7750
rect 16120 7686 16172 7692
rect 16132 6322 16160 7686
rect 16316 7002 16344 7754
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16592 6458 16620 8366
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16684 6390 16712 8298
rect 16776 7546 16804 11494
rect 17144 11218 17172 12702
rect 17222 12744 17278 12753
rect 17222 12679 17278 12688
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16672 6384 16724 6390
rect 16672 6326 16724 6332
rect 16776 6322 16804 7482
rect 16960 7290 16988 10950
rect 17236 10606 17264 12679
rect 17328 10810 17356 13262
rect 17972 13258 18000 14878
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 18064 13870 18092 14214
rect 18156 14074 18184 15370
rect 18248 14074 18276 16390
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18524 14006 18552 16934
rect 18604 16516 18656 16522
rect 18604 16458 18656 16464
rect 18616 14482 18644 16458
rect 18892 15638 18920 17750
rect 19352 17678 19380 19314
rect 19536 18222 19564 19382
rect 19616 19236 19668 19242
rect 19616 19178 19668 19184
rect 19628 18222 19656 19178
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19720 18358 19748 19110
rect 19812 18698 19840 20198
rect 19916 20156 20292 20165
rect 19972 20154 19996 20156
rect 20052 20154 20076 20156
rect 20132 20154 20156 20156
rect 20212 20154 20236 20156
rect 19972 20102 19982 20154
rect 20226 20102 20236 20154
rect 19972 20100 19996 20102
rect 20052 20100 20076 20102
rect 20132 20100 20156 20102
rect 20212 20100 20236 20102
rect 19916 20091 20292 20100
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 20656 19612 21032 19621
rect 20712 19610 20736 19612
rect 20792 19610 20816 19612
rect 20872 19610 20896 19612
rect 20952 19610 20976 19612
rect 20712 19558 20722 19610
rect 20966 19558 20976 19610
rect 20712 19556 20736 19558
rect 20792 19556 20816 19558
rect 20872 19556 20896 19558
rect 20952 19556 20976 19558
rect 20656 19547 21032 19556
rect 21376 19514 21404 19654
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 20444 19304 20496 19310
rect 20444 19246 20496 19252
rect 19916 19068 20292 19077
rect 19972 19066 19996 19068
rect 20052 19066 20076 19068
rect 20132 19066 20156 19068
rect 20212 19066 20236 19068
rect 19972 19014 19982 19066
rect 20226 19014 20236 19066
rect 19972 19012 19996 19014
rect 20052 19012 20076 19014
rect 20132 19012 20156 19014
rect 20212 19012 20236 19014
rect 19916 19003 20292 19012
rect 20456 18970 20484 19246
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 21468 18766 21496 20198
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23308 19145 23336 19314
rect 23294 19136 23350 19145
rect 23294 19071 23350 19080
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 19800 18692 19852 18698
rect 19800 18634 19852 18640
rect 20656 18524 21032 18533
rect 20712 18522 20736 18524
rect 20792 18522 20816 18524
rect 20872 18522 20896 18524
rect 20952 18522 20976 18524
rect 20712 18470 20722 18522
rect 20966 18470 20976 18522
rect 20712 18468 20736 18470
rect 20792 18468 20816 18470
rect 20872 18468 20896 18470
rect 20952 18468 20976 18470
rect 20656 18459 21032 18468
rect 21284 18426 21312 18702
rect 23296 18692 23348 18698
rect 23296 18634 23348 18640
rect 23308 18465 23336 18634
rect 23294 18456 23350 18465
rect 21272 18420 21324 18426
rect 23294 18391 23350 18400
rect 21272 18362 21324 18368
rect 19708 18352 19760 18358
rect 19708 18294 19760 18300
rect 19524 18216 19576 18222
rect 19524 18158 19576 18164
rect 19616 18216 19668 18222
rect 19616 18158 19668 18164
rect 19064 17672 19116 17678
rect 19064 17614 19116 17620
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18984 17338 19012 17478
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 19076 15978 19104 17614
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19248 16448 19300 16454
rect 19248 16390 19300 16396
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19064 15972 19116 15978
rect 19064 15914 19116 15920
rect 18880 15632 18932 15638
rect 18880 15574 18932 15580
rect 19260 15094 19288 16390
rect 19352 15706 19380 16390
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 19444 15026 19472 17478
rect 19536 16998 19564 18158
rect 19916 17980 20292 17989
rect 19972 17978 19996 17980
rect 20052 17978 20076 17980
rect 20132 17978 20156 17980
rect 20212 17978 20236 17980
rect 19972 17926 19982 17978
rect 20226 17926 20236 17978
rect 19972 17924 19996 17926
rect 20052 17924 20076 17926
rect 20132 17924 20156 17926
rect 20212 17924 20236 17926
rect 19916 17915 20292 17924
rect 20656 17436 21032 17445
rect 20712 17434 20736 17436
rect 20792 17434 20816 17436
rect 20872 17434 20896 17436
rect 20952 17434 20976 17436
rect 20712 17382 20722 17434
rect 20966 17382 20976 17434
rect 20712 17380 20736 17382
rect 20792 17380 20816 17382
rect 20872 17380 20896 17382
rect 20952 17380 20976 17382
rect 20656 17371 21032 17380
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 21180 17196 21232 17202
rect 21180 17138 21232 17144
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19536 16250 19564 16934
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 19524 15428 19576 15434
rect 19524 15370 19576 15376
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19536 14958 19564 15370
rect 19628 15366 19656 17138
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 19916 16892 20292 16901
rect 19972 16890 19996 16892
rect 20052 16890 20076 16892
rect 20132 16890 20156 16892
rect 20212 16890 20236 16892
rect 19972 16838 19982 16890
rect 20226 16838 20236 16890
rect 19972 16836 19996 16838
rect 20052 16836 20076 16838
rect 20132 16836 20156 16838
rect 20212 16836 20236 16838
rect 19916 16827 20292 16836
rect 19892 16788 19944 16794
rect 19892 16730 19944 16736
rect 19800 16720 19852 16726
rect 19800 16662 19852 16668
rect 19708 16448 19760 16454
rect 19708 16390 19760 16396
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19720 15094 19748 16390
rect 19812 16250 19840 16662
rect 19800 16244 19852 16250
rect 19800 16186 19852 16192
rect 19904 15994 19932 16730
rect 21100 16658 21128 16934
rect 21192 16794 21220 17138
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 21732 16720 21784 16726
rect 21732 16662 21784 16668
rect 21088 16652 21140 16658
rect 21088 16594 21140 16600
rect 20656 16348 21032 16357
rect 20712 16346 20736 16348
rect 20792 16346 20816 16348
rect 20872 16346 20896 16348
rect 20952 16346 20976 16348
rect 20712 16294 20722 16346
rect 20966 16294 20976 16346
rect 20712 16292 20736 16294
rect 20792 16292 20816 16294
rect 20872 16292 20896 16294
rect 20952 16292 20976 16294
rect 20656 16283 21032 16292
rect 19812 15966 19932 15994
rect 20352 16040 20404 16046
rect 20352 15982 20404 15988
rect 19708 15088 19760 15094
rect 19708 15030 19760 15036
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19812 14822 19840 15966
rect 19916 15804 20292 15813
rect 19972 15802 19996 15804
rect 20052 15802 20076 15804
rect 20132 15802 20156 15804
rect 20212 15802 20236 15804
rect 19972 15750 19982 15802
rect 20226 15750 20236 15802
rect 19972 15748 19996 15750
rect 20052 15748 20076 15750
rect 20132 15748 20156 15750
rect 20212 15748 20236 15750
rect 19916 15739 20292 15748
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19916 14716 20292 14725
rect 19972 14714 19996 14716
rect 20052 14714 20076 14716
rect 20132 14714 20156 14716
rect 20212 14714 20236 14716
rect 19972 14662 19982 14714
rect 20226 14662 20236 14714
rect 19972 14660 19996 14662
rect 20052 14660 20076 14662
rect 20132 14660 20156 14662
rect 20212 14660 20236 14662
rect 19916 14651 20292 14660
rect 20364 14600 20392 15982
rect 21640 15972 21692 15978
rect 21640 15914 21692 15920
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21088 15632 21140 15638
rect 21088 15574 21140 15580
rect 20656 15260 21032 15269
rect 20712 15258 20736 15260
rect 20792 15258 20816 15260
rect 20872 15258 20896 15260
rect 20952 15258 20976 15260
rect 20712 15206 20722 15258
rect 20966 15206 20976 15258
rect 20712 15204 20736 15206
rect 20792 15204 20816 15206
rect 20872 15204 20896 15206
rect 20952 15204 20976 15206
rect 20656 15195 21032 15204
rect 21100 15162 21128 15574
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20548 14618 20576 14758
rect 20088 14572 20392 14600
rect 20536 14612 20588 14618
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18616 14278 18644 14418
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19800 14340 19852 14346
rect 19800 14282 19852 14288
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18972 14272 19024 14278
rect 18972 14214 19024 14220
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18052 13320 18104 13326
rect 18104 13280 18276 13308
rect 18052 13262 18104 13268
rect 17960 13252 18012 13258
rect 17960 13194 18012 13200
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17604 12306 17632 12582
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17512 10810 17540 12242
rect 17592 11620 17644 11626
rect 17592 11562 17644 11568
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17604 9994 17632 11562
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17788 10266 17816 10950
rect 17972 10742 18000 13194
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18156 12374 18184 13126
rect 18144 12368 18196 12374
rect 18144 12310 18196 12316
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 18156 9994 18184 12174
rect 18248 9994 18276 13280
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18892 12986 18920 13126
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 18984 12434 19012 14214
rect 19352 14074 19380 14282
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19260 12986 19288 13126
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 18984 12406 19104 12434
rect 19076 12238 19104 12406
rect 19064 12232 19116 12238
rect 19064 12174 19116 12180
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18432 10742 18460 12038
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18512 11212 18564 11218
rect 18512 11154 18564 11160
rect 18420 10736 18472 10742
rect 18420 10678 18472 10684
rect 18524 9994 18552 11154
rect 17592 9988 17644 9994
rect 17592 9930 17644 9936
rect 18144 9988 18196 9994
rect 18144 9930 18196 9936
rect 18236 9988 18288 9994
rect 18236 9930 18288 9936
rect 18512 9988 18564 9994
rect 18512 9930 18564 9936
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 17144 8498 17172 9862
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17420 9178 17448 9318
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17604 9042 17632 9930
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17684 7812 17736 7818
rect 17684 7754 17736 7760
rect 16960 7262 17172 7290
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 16684 4826 16712 5646
rect 16960 5234 16988 7142
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14656 4380 15032 4389
rect 14712 4378 14736 4380
rect 14792 4378 14816 4380
rect 14872 4378 14896 4380
rect 14952 4378 14976 4380
rect 14712 4326 14722 4378
rect 14966 4326 14976 4378
rect 14712 4324 14736 4326
rect 14792 4324 14816 4326
rect 14872 4324 14896 4326
rect 14952 4324 14976 4326
rect 14656 4315 15032 4324
rect 14372 4004 14424 4010
rect 14372 3946 14424 3952
rect 13916 3836 14292 3845
rect 13972 3834 13996 3836
rect 14052 3834 14076 3836
rect 14132 3834 14156 3836
rect 14212 3834 14236 3836
rect 13972 3782 13982 3834
rect 14226 3782 14236 3834
rect 13972 3780 13996 3782
rect 14052 3780 14076 3782
rect 14132 3780 14156 3782
rect 14212 3780 14236 3782
rect 13916 3771 14292 3780
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 14656 3292 15032 3301
rect 14712 3290 14736 3292
rect 14792 3290 14816 3292
rect 14872 3290 14896 3292
rect 14952 3290 14976 3292
rect 14712 3238 14722 3290
rect 14966 3238 14976 3290
rect 14712 3236 14736 3238
rect 14792 3236 14816 3238
rect 14872 3236 14896 3238
rect 14952 3236 14976 3238
rect 14656 3227 15032 3236
rect 13916 2748 14292 2757
rect 13972 2746 13996 2748
rect 14052 2746 14076 2748
rect 14132 2746 14156 2748
rect 14212 2746 14236 2748
rect 13972 2694 13982 2746
rect 14226 2694 14236 2746
rect 13972 2692 13996 2694
rect 14052 2692 14076 2694
rect 14132 2692 14156 2694
rect 14212 2692 14236 2694
rect 13916 2683 14292 2692
rect 17052 2446 17080 6054
rect 17144 4826 17172 7262
rect 17696 6662 17724 7754
rect 17880 6730 17908 9386
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17972 8906 18000 9318
rect 18524 8906 18552 9930
rect 18616 9110 18644 11698
rect 18972 10736 19024 10742
rect 18972 10678 19024 10684
rect 18880 10192 18932 10198
rect 18880 10134 18932 10140
rect 18604 9104 18656 9110
rect 18604 9046 18656 9052
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 18512 8900 18564 8906
rect 18512 8842 18564 8848
rect 18696 8900 18748 8906
rect 18696 8842 18748 8848
rect 17972 8498 18000 8842
rect 18524 8566 18552 8842
rect 18512 8560 18564 8566
rect 18512 8502 18564 8508
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17696 5778 17724 6598
rect 18064 5914 18092 7278
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18156 5846 18184 6258
rect 18144 5840 18196 5846
rect 18144 5782 18196 5788
rect 17684 5772 17736 5778
rect 17684 5714 17736 5720
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17420 5370 17448 5578
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 18064 2774 18092 5510
rect 18248 5234 18276 8298
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18340 5710 18368 7346
rect 18524 6458 18552 7754
rect 18708 7750 18736 8842
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18800 6458 18828 8774
rect 18892 8430 18920 10134
rect 18880 8424 18932 8430
rect 18880 8366 18932 8372
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18892 7002 18920 7822
rect 18880 6996 18932 7002
rect 18880 6938 18932 6944
rect 18984 6798 19012 10678
rect 19352 10554 19380 13262
rect 19812 12986 19840 14282
rect 20088 13954 20116 14572
rect 20536 14554 20588 14560
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 19996 13938 20116 13954
rect 19984 13932 20116 13938
rect 20036 13926 20116 13932
rect 19984 13874 20036 13880
rect 19916 13628 20292 13637
rect 19972 13626 19996 13628
rect 20052 13626 20076 13628
rect 20132 13626 20156 13628
rect 20212 13626 20236 13628
rect 19972 13574 19982 13626
rect 20226 13574 20236 13626
rect 19972 13572 19996 13574
rect 20052 13572 20076 13574
rect 20132 13572 20156 13574
rect 20212 13572 20236 13574
rect 19916 13563 20292 13572
rect 19892 13524 19944 13530
rect 19892 13466 19944 13472
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 19904 12850 19932 13466
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19616 12844 19668 12850
rect 19616 12786 19668 12792
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19628 11014 19656 12786
rect 19996 12782 20024 13126
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 20456 12646 20484 14350
rect 20640 14278 20668 14894
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 20656 14172 21032 14181
rect 20712 14170 20736 14172
rect 20792 14170 20816 14172
rect 20872 14170 20896 14172
rect 20952 14170 20976 14172
rect 20712 14118 20722 14170
rect 20966 14118 20976 14170
rect 20712 14116 20736 14118
rect 20792 14116 20816 14118
rect 20872 14116 20896 14118
rect 20952 14116 20976 14118
rect 20656 14107 21032 14116
rect 20812 13728 20864 13734
rect 20812 13670 20864 13676
rect 20824 13258 20852 13670
rect 20812 13252 20864 13258
rect 20812 13194 20864 13200
rect 20656 13084 21032 13093
rect 20712 13082 20736 13084
rect 20792 13082 20816 13084
rect 20872 13082 20896 13084
rect 20952 13082 20976 13084
rect 20712 13030 20722 13082
rect 20966 13030 20976 13082
rect 20712 13028 20736 13030
rect 20792 13028 20816 13030
rect 20872 13028 20896 13030
rect 20952 13028 20976 13030
rect 20656 13019 21032 13028
rect 21100 12850 21128 15098
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21192 13870 21220 14214
rect 21284 14074 21312 14758
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21376 13870 21404 15302
rect 21468 13938 21496 15846
rect 21652 15094 21680 15914
rect 21640 15088 21692 15094
rect 21640 15030 21692 15036
rect 21744 13938 21772 16662
rect 22192 16652 22244 16658
rect 22192 16594 22244 16600
rect 21916 16448 21968 16454
rect 21916 16390 21968 16396
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 21548 13932 21600 13938
rect 21548 13874 21600 13880
rect 21732 13932 21784 13938
rect 21732 13874 21784 13880
rect 21180 13864 21232 13870
rect 21180 13806 21232 13812
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21560 13433 21588 13874
rect 21546 13424 21602 13433
rect 21546 13359 21602 13368
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 21364 12844 21416 12850
rect 21364 12786 21416 12792
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 19916 12540 20292 12549
rect 19972 12538 19996 12540
rect 20052 12538 20076 12540
rect 20132 12538 20156 12540
rect 20212 12538 20236 12540
rect 19972 12486 19982 12538
rect 20226 12486 20236 12538
rect 19972 12484 19996 12486
rect 20052 12484 20076 12486
rect 20132 12484 20156 12486
rect 20212 12484 20236 12486
rect 19916 12475 20292 12484
rect 21180 12300 21232 12306
rect 21180 12242 21232 12248
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19720 11218 19748 12174
rect 20444 12164 20496 12170
rect 20444 12106 20496 12112
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19076 10538 19380 10554
rect 19064 10532 19380 10538
rect 19116 10526 19380 10532
rect 19064 10474 19116 10480
rect 19156 10464 19208 10470
rect 19156 10406 19208 10412
rect 19168 9994 19196 10406
rect 19444 10282 19472 10610
rect 19812 10577 19840 11494
rect 19916 11452 20292 11461
rect 19972 11450 19996 11452
rect 20052 11450 20076 11452
rect 20132 11450 20156 11452
rect 20212 11450 20236 11452
rect 19972 11398 19982 11450
rect 20226 11398 20236 11450
rect 19972 11396 19996 11398
rect 20052 11396 20076 11398
rect 20132 11396 20156 11398
rect 20212 11396 20236 11398
rect 19916 11387 20292 11396
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 19798 10568 19854 10577
rect 19798 10503 19854 10512
rect 19916 10364 20292 10373
rect 19972 10362 19996 10364
rect 20052 10362 20076 10364
rect 20132 10362 20156 10364
rect 20212 10362 20236 10364
rect 19972 10310 19982 10362
rect 20226 10310 20236 10362
rect 19972 10308 19996 10310
rect 20052 10308 20076 10310
rect 20132 10308 20156 10310
rect 20212 10308 20236 10310
rect 19916 10299 20292 10308
rect 19352 10254 19472 10282
rect 20364 10266 20392 11086
rect 20456 10674 20484 12106
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 20548 11830 20576 12038
rect 20656 11996 21032 12005
rect 20712 11994 20736 11996
rect 20792 11994 20816 11996
rect 20872 11994 20896 11996
rect 20952 11994 20976 11996
rect 20712 11942 20722 11994
rect 20966 11942 20976 11994
rect 20712 11940 20736 11942
rect 20792 11940 20816 11942
rect 20872 11940 20896 11942
rect 20952 11940 20976 11942
rect 20656 11931 21032 11940
rect 21100 11898 21128 12038
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 20536 11824 20588 11830
rect 20536 11766 20588 11772
rect 21192 11558 21220 12242
rect 21376 11830 21404 12786
rect 21560 11898 21588 13262
rect 21640 12912 21692 12918
rect 21640 12854 21692 12860
rect 21652 11898 21680 12854
rect 21744 12782 21772 13874
rect 21824 13320 21876 13326
rect 21824 13262 21876 13268
rect 21732 12776 21784 12782
rect 21732 12718 21784 12724
rect 21732 12640 21784 12646
rect 21732 12582 21784 12588
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 21364 11824 21416 11830
rect 21364 11766 21416 11772
rect 21640 11756 21692 11762
rect 21640 11698 21692 11704
rect 21180 11552 21232 11558
rect 21180 11494 21232 11500
rect 21086 11248 21142 11257
rect 21086 11183 21142 11192
rect 21548 11212 21600 11218
rect 20656 10908 21032 10917
rect 20712 10906 20736 10908
rect 20792 10906 20816 10908
rect 20872 10906 20896 10908
rect 20952 10906 20976 10908
rect 20712 10854 20722 10906
rect 20966 10854 20976 10906
rect 20712 10852 20736 10854
rect 20792 10852 20816 10854
rect 20872 10852 20896 10854
rect 20952 10852 20976 10854
rect 20656 10843 21032 10852
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 20904 10600 20956 10606
rect 20904 10542 20956 10548
rect 19352 10062 19380 10254
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19156 9988 19208 9994
rect 19156 9930 19208 9936
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 18788 6452 18840 6458
rect 18788 6394 18840 6400
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18340 5234 18368 5646
rect 18432 5370 18460 6190
rect 18420 5364 18472 5370
rect 18420 5306 18472 5312
rect 19076 5234 19104 8570
rect 19168 5710 19196 9114
rect 19248 9104 19300 9110
rect 19300 9052 19380 9058
rect 19248 9046 19380 9052
rect 19260 9030 19380 9046
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19260 6458 19288 6734
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19352 5778 19380 9030
rect 19444 7410 19472 10254
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19444 7002 19472 7346
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19536 6882 19564 9590
rect 20088 9489 20116 9998
rect 20916 9926 20944 10542
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 20656 9820 21032 9829
rect 20712 9818 20736 9820
rect 20792 9818 20816 9820
rect 20872 9818 20896 9820
rect 20952 9818 20976 9820
rect 20712 9766 20722 9818
rect 20966 9766 20976 9818
rect 20712 9764 20736 9766
rect 20792 9764 20816 9766
rect 20872 9764 20896 9766
rect 20952 9764 20976 9766
rect 20656 9755 21032 9764
rect 21100 9674 21128 11183
rect 21548 11154 21600 11160
rect 21456 11008 21508 11014
rect 21456 10950 21508 10956
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 21178 10296 21234 10305
rect 21178 10231 21234 10240
rect 21008 9646 21128 9674
rect 20810 9616 20866 9625
rect 20810 9551 20812 9560
rect 20864 9551 20866 9560
rect 20812 9522 20864 9528
rect 20074 9480 20130 9489
rect 20074 9415 20130 9424
rect 20352 9444 20404 9450
rect 20352 9386 20404 9392
rect 19916 9276 20292 9285
rect 19972 9274 19996 9276
rect 20052 9274 20076 9276
rect 20132 9274 20156 9276
rect 20212 9274 20236 9276
rect 19972 9222 19982 9274
rect 20226 9222 20236 9274
rect 19972 9220 19996 9222
rect 20052 9220 20076 9222
rect 20132 9220 20156 9222
rect 20212 9220 20236 9222
rect 19916 9211 20292 9220
rect 20364 9110 20392 9386
rect 20352 9104 20404 9110
rect 20352 9046 20404 9052
rect 20536 9104 20588 9110
rect 20536 9046 20588 9052
rect 20548 8566 20576 9046
rect 21008 8820 21036 9646
rect 21192 9625 21220 10231
rect 21270 10160 21326 10169
rect 21270 10095 21326 10104
rect 21178 9616 21234 9625
rect 21178 9551 21234 9560
rect 21008 8792 21128 8820
rect 20656 8732 21032 8741
rect 20712 8730 20736 8732
rect 20792 8730 20816 8732
rect 20872 8730 20896 8732
rect 20952 8730 20976 8732
rect 20712 8678 20722 8730
rect 20966 8678 20976 8730
rect 20712 8676 20736 8678
rect 20792 8676 20816 8678
rect 20872 8676 20896 8678
rect 20952 8676 20976 8678
rect 20656 8667 21032 8676
rect 20536 8560 20588 8566
rect 20536 8502 20588 8508
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19444 6854 19564 6882
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19156 5704 19208 5710
rect 19156 5646 19208 5652
rect 19168 5370 19196 5646
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 19064 5228 19116 5234
rect 19064 5170 19116 5176
rect 19076 4622 19104 5170
rect 19444 5166 19472 6854
rect 19524 6724 19576 6730
rect 19524 6666 19576 6672
rect 19536 5846 19564 6666
rect 19628 5914 19656 7278
rect 19720 6730 19748 7346
rect 19708 6724 19760 6730
rect 19708 6666 19760 6672
rect 19812 6322 19840 8366
rect 19916 8188 20292 8197
rect 19972 8186 19996 8188
rect 20052 8186 20076 8188
rect 20132 8186 20156 8188
rect 20212 8186 20236 8188
rect 19972 8134 19982 8186
rect 20226 8134 20236 8186
rect 19972 8132 19996 8134
rect 20052 8132 20076 8134
rect 20132 8132 20156 8134
rect 20212 8132 20236 8134
rect 19916 8123 20292 8132
rect 19916 7100 20292 7109
rect 19972 7098 19996 7100
rect 20052 7098 20076 7100
rect 20132 7098 20156 7100
rect 20212 7098 20236 7100
rect 19972 7046 19982 7098
rect 20226 7046 20236 7098
rect 19972 7044 19996 7046
rect 20052 7044 20076 7046
rect 20132 7044 20156 7046
rect 20212 7044 20236 7046
rect 19916 7035 20292 7044
rect 19800 6316 19852 6322
rect 19800 6258 19852 6264
rect 20352 6112 20404 6118
rect 20352 6054 20404 6060
rect 19916 6012 20292 6021
rect 19972 6010 19996 6012
rect 20052 6010 20076 6012
rect 20132 6010 20156 6012
rect 20212 6010 20236 6012
rect 19972 5958 19982 6010
rect 20226 5958 20236 6010
rect 19972 5956 19996 5958
rect 20052 5956 20076 5958
rect 20132 5956 20156 5958
rect 20212 5956 20236 5958
rect 19916 5947 20292 5956
rect 20364 5914 20392 6054
rect 19616 5908 19668 5914
rect 19616 5850 19668 5856
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 19524 5840 19576 5846
rect 20456 5794 20484 8434
rect 20656 7644 21032 7653
rect 20712 7642 20736 7644
rect 20792 7642 20816 7644
rect 20872 7642 20896 7644
rect 20952 7642 20976 7644
rect 20712 7590 20722 7642
rect 20966 7590 20976 7642
rect 20712 7588 20736 7590
rect 20792 7588 20816 7590
rect 20872 7588 20896 7590
rect 20952 7588 20976 7590
rect 20656 7579 21032 7588
rect 21100 7546 21128 8792
rect 21192 8294 21220 9551
rect 21284 8634 21312 10095
rect 21376 9722 21404 10610
rect 21468 10305 21496 10950
rect 21454 10296 21510 10305
rect 21454 10231 21510 10240
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21364 9512 21416 9518
rect 21362 9480 21364 9489
rect 21416 9480 21418 9489
rect 21362 9415 21418 9424
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21180 7744 21232 7750
rect 21180 7686 21232 7692
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 20656 6556 21032 6565
rect 20712 6554 20736 6556
rect 20792 6554 20816 6556
rect 20872 6554 20896 6556
rect 20952 6554 20976 6556
rect 20712 6502 20722 6554
rect 20966 6502 20976 6554
rect 20712 6500 20736 6502
rect 20792 6500 20816 6502
rect 20872 6500 20896 6502
rect 20952 6500 20976 6502
rect 20656 6491 21032 6500
rect 20996 6384 21048 6390
rect 20996 6326 21048 6332
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20916 5914 20944 6054
rect 21008 5914 21036 6326
rect 21192 6322 21220 7686
rect 21284 7546 21312 8570
rect 21376 8090 21404 8910
rect 21364 8084 21416 8090
rect 21364 8026 21416 8032
rect 21468 7546 21496 9998
rect 21560 8480 21588 11154
rect 21652 10606 21680 11698
rect 21640 10600 21692 10606
rect 21640 10542 21692 10548
rect 21640 9920 21692 9926
rect 21640 9862 21692 9868
rect 21652 9489 21680 9862
rect 21744 9625 21772 12582
rect 21836 12306 21864 13262
rect 21824 12300 21876 12306
rect 21824 12242 21876 12248
rect 21928 11762 21956 16390
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 21916 11756 21968 11762
rect 21916 11698 21968 11704
rect 21824 11688 21876 11694
rect 21824 11630 21876 11636
rect 21730 9616 21786 9625
rect 21730 9551 21786 9560
rect 21744 9518 21772 9551
rect 21732 9512 21784 9518
rect 21638 9480 21694 9489
rect 21732 9454 21784 9460
rect 21638 9415 21694 9424
rect 21744 8498 21772 9454
rect 21836 8634 21864 11630
rect 22020 11286 22048 16050
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 22112 15162 22140 15982
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 22112 14074 22140 14350
rect 22100 14068 22152 14074
rect 22100 14010 22152 14016
rect 22204 13530 22232 16594
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22572 15502 22600 15846
rect 22560 15496 22612 15502
rect 22560 15438 22612 15444
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22560 15360 22612 15366
rect 22560 15302 22612 15308
rect 22376 15020 22428 15026
rect 22376 14962 22428 14968
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22296 14414 22324 14758
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22204 12918 22232 13466
rect 22388 13326 22416 14962
rect 22468 14816 22520 14822
rect 22468 14758 22520 14764
rect 22376 13320 22428 13326
rect 22376 13262 22428 13268
rect 22192 12912 22244 12918
rect 22192 12854 22244 12860
rect 22376 12844 22428 12850
rect 22296 12804 22376 12832
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 22100 11076 22152 11082
rect 22100 11018 22152 11024
rect 22008 11008 22060 11014
rect 22008 10950 22060 10956
rect 21916 10668 21968 10674
rect 21916 10610 21968 10616
rect 21928 9994 21956 10610
rect 22020 10062 22048 10950
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 21916 9988 21968 9994
rect 21916 9930 21968 9936
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21640 8492 21692 8498
rect 21560 8452 21640 8480
rect 21640 8434 21692 8440
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 21652 7886 21680 8434
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 21548 7880 21600 7886
rect 21548 7822 21600 7828
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21284 6322 21312 7482
rect 21456 7268 21508 7274
rect 21456 7210 21508 7216
rect 21364 6792 21416 6798
rect 21364 6734 21416 6740
rect 21180 6316 21232 6322
rect 21180 6258 21232 6264
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 19524 5782 19576 5788
rect 20180 5766 20484 5794
rect 20180 5710 20208 5766
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 21272 5636 21324 5642
rect 21272 5578 21324 5584
rect 20656 5468 21032 5477
rect 20712 5466 20736 5468
rect 20792 5466 20816 5468
rect 20872 5466 20896 5468
rect 20952 5466 20976 5468
rect 20712 5414 20722 5466
rect 20966 5414 20976 5466
rect 20712 5412 20736 5414
rect 20792 5412 20816 5414
rect 20872 5412 20896 5414
rect 20952 5412 20976 5414
rect 20656 5403 21032 5412
rect 21284 5370 21312 5578
rect 21376 5370 21404 6734
rect 21468 5778 21496 7210
rect 21560 5914 21588 7822
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 21456 5772 21508 5778
rect 21456 5714 21508 5720
rect 21652 5642 21680 7822
rect 21732 7812 21784 7818
rect 21732 7754 21784 7760
rect 21640 5636 21692 5642
rect 21640 5578 21692 5584
rect 21272 5364 21324 5370
rect 21272 5306 21324 5312
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19916 4924 20292 4933
rect 19972 4922 19996 4924
rect 20052 4922 20076 4924
rect 20132 4922 20156 4924
rect 20212 4922 20236 4924
rect 19972 4870 19982 4922
rect 20226 4870 20236 4922
rect 19972 4868 19996 4870
rect 20052 4868 20076 4870
rect 20132 4868 20156 4870
rect 20212 4868 20236 4870
rect 19916 4859 20292 4868
rect 21744 4826 21772 7754
rect 21836 5778 21864 7890
rect 21928 7410 21956 9522
rect 22112 8922 22140 11018
rect 22296 10169 22324 12804
rect 22376 12786 22428 12792
rect 22480 11558 22508 14758
rect 22572 14346 22600 15302
rect 22664 14618 22692 15438
rect 22652 14612 22704 14618
rect 22652 14554 22704 14560
rect 22560 14340 22612 14346
rect 22560 14282 22612 14288
rect 22664 14006 22692 14554
rect 22652 14000 22704 14006
rect 22652 13942 22704 13948
rect 22560 12640 22612 12646
rect 22560 12582 22612 12588
rect 22572 11830 22600 12582
rect 22650 12336 22706 12345
rect 22650 12271 22706 12280
rect 22560 11824 22612 11830
rect 22560 11766 22612 11772
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22466 10976 22522 10985
rect 22466 10911 22522 10920
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22282 10160 22338 10169
rect 22282 10095 22338 10104
rect 22112 8894 22324 8922
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 22008 6996 22060 7002
rect 22008 6938 22060 6944
rect 22020 5914 22048 6938
rect 22008 5908 22060 5914
rect 22008 5850 22060 5856
rect 21824 5772 21876 5778
rect 21824 5714 21876 5720
rect 21732 4820 21784 4826
rect 21732 4762 21784 4768
rect 22112 4690 22140 8774
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 22204 6866 22232 8570
rect 22296 7002 22324 8894
rect 22284 6996 22336 7002
rect 22284 6938 22336 6944
rect 22192 6860 22244 6866
rect 22192 6802 22244 6808
rect 22388 5370 22416 10746
rect 22480 10062 22508 10911
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22664 9042 22692 12271
rect 22756 10656 22784 16390
rect 22928 16040 22980 16046
rect 22928 15982 22980 15988
rect 22836 15904 22888 15910
rect 22836 15846 22888 15852
rect 22848 14226 22876 15846
rect 22940 14362 22968 15982
rect 23032 15434 23060 16526
rect 23204 16516 23256 16522
rect 23204 16458 23256 16464
rect 23112 16448 23164 16454
rect 23112 16390 23164 16396
rect 23124 16182 23152 16390
rect 23112 16176 23164 16182
rect 23112 16118 23164 16124
rect 23216 16130 23244 16458
rect 23308 16425 23336 17070
rect 23294 16416 23350 16425
rect 23294 16351 23350 16360
rect 23020 15428 23072 15434
rect 23020 15370 23072 15376
rect 23124 15366 23152 16118
rect 23216 16102 23336 16130
rect 23204 15972 23256 15978
rect 23204 15914 23256 15920
rect 23112 15360 23164 15366
rect 23112 15302 23164 15308
rect 22940 14334 23060 14362
rect 22848 14198 22968 14226
rect 22836 12776 22888 12782
rect 22836 12718 22888 12724
rect 22848 12102 22876 12718
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 22940 10810 22968 14198
rect 23032 11626 23060 14334
rect 23124 12442 23152 15302
rect 23216 15026 23244 15914
rect 23308 15745 23336 16102
rect 23294 15736 23350 15745
rect 23294 15671 23350 15680
rect 23204 15020 23256 15026
rect 23204 14962 23256 14968
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 23204 14884 23256 14890
rect 23204 14826 23256 14832
rect 23216 14006 23244 14826
rect 23308 14006 23336 14962
rect 23386 14376 23442 14385
rect 23386 14311 23388 14320
rect 23440 14311 23442 14320
rect 23388 14282 23440 14288
rect 23204 14000 23256 14006
rect 23204 13942 23256 13948
rect 23296 14000 23348 14006
rect 23296 13942 23348 13948
rect 23386 13696 23442 13705
rect 23386 13631 23442 13640
rect 23400 13394 23428 13631
rect 23388 13388 23440 13394
rect 23388 13330 23440 13336
rect 23388 13252 23440 13258
rect 23388 13194 23440 13200
rect 23400 13025 23428 13194
rect 23386 13016 23442 13025
rect 23386 12951 23442 12960
rect 23112 12436 23164 12442
rect 23112 12378 23164 12384
rect 23388 12436 23440 12442
rect 23388 12378 23440 12384
rect 23296 11756 23348 11762
rect 23296 11698 23348 11704
rect 23202 11656 23258 11665
rect 23020 11620 23072 11626
rect 23202 11591 23258 11600
rect 23020 11562 23072 11568
rect 23110 11248 23166 11257
rect 23110 11183 23166 11192
rect 23124 11150 23152 11183
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 23112 11144 23164 11150
rect 23112 11086 23164 11092
rect 23032 10810 23060 11086
rect 23216 10826 23244 11591
rect 23308 11354 23336 11698
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 22928 10804 22980 10810
rect 22928 10746 22980 10752
rect 23020 10804 23072 10810
rect 23216 10798 23336 10826
rect 23020 10746 23072 10752
rect 23204 10668 23256 10674
rect 22756 10628 23204 10656
rect 23204 10610 23256 10616
rect 22742 10568 22798 10577
rect 22742 10503 22798 10512
rect 22756 10062 22784 10503
rect 23308 10130 23336 10798
rect 23296 10124 23348 10130
rect 23296 10066 23348 10072
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 23294 9480 23350 9489
rect 23294 9415 23296 9424
rect 23348 9415 23350 9424
rect 23296 9386 23348 9392
rect 23112 9376 23164 9382
rect 23112 9318 23164 9324
rect 22652 9036 22704 9042
rect 22652 8978 22704 8984
rect 23018 8936 23074 8945
rect 22940 8894 23018 8922
rect 22468 8288 22520 8294
rect 22468 8230 22520 8236
rect 22376 5364 22428 5370
rect 22376 5306 22428 5312
rect 22480 5234 22508 8230
rect 22744 7812 22796 7818
rect 22744 7754 22796 7760
rect 22560 6656 22612 6662
rect 22560 6598 22612 6604
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 22100 4684 22152 4690
rect 22100 4626 22152 4632
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 20656 4380 21032 4389
rect 20712 4378 20736 4380
rect 20792 4378 20816 4380
rect 20872 4378 20896 4380
rect 20952 4378 20976 4380
rect 20712 4326 20722 4378
rect 20966 4326 20976 4378
rect 20712 4324 20736 4326
rect 20792 4324 20816 4326
rect 20872 4324 20896 4326
rect 20952 4324 20976 4326
rect 20656 4315 21032 4324
rect 22572 4146 22600 6598
rect 22756 4826 22784 7754
rect 22940 6866 22968 8894
rect 23018 8871 23074 8880
rect 23020 7880 23072 7886
rect 23020 7822 23072 7828
rect 22928 6860 22980 6866
rect 22928 6802 22980 6808
rect 23032 6458 23060 7822
rect 23124 7410 23152 9318
rect 23296 8832 23348 8838
rect 23296 8774 23348 8780
rect 23308 8498 23336 8774
rect 23296 8492 23348 8498
rect 23296 8434 23348 8440
rect 23294 8256 23350 8265
rect 23216 8214 23294 8242
rect 23112 7404 23164 7410
rect 23112 7346 23164 7352
rect 23216 6882 23244 8214
rect 23294 8191 23350 8200
rect 23296 7880 23348 7886
rect 23296 7822 23348 7828
rect 23308 7478 23336 7822
rect 23296 7472 23348 7478
rect 23296 7414 23348 7420
rect 23216 6854 23336 6882
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 22744 4820 22796 4826
rect 22744 4762 22796 4768
rect 23124 4146 23152 6258
rect 23204 6248 23256 6254
rect 23204 6190 23256 6196
rect 23216 5370 23244 6190
rect 23308 5710 23336 6854
rect 23400 6322 23428 12378
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 23492 9586 23520 12174
rect 23480 9580 23532 9586
rect 23480 9522 23532 9528
rect 23480 7200 23532 7206
rect 23480 7142 23532 7148
rect 23388 6316 23440 6322
rect 23388 6258 23440 6264
rect 23400 5710 23428 6258
rect 23296 5704 23348 5710
rect 23296 5646 23348 5652
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 23204 5364 23256 5370
rect 23204 5306 23256 5312
rect 23400 5234 23428 5646
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 23492 4690 23520 7142
rect 23480 4684 23532 4690
rect 23480 4626 23532 4632
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 19916 3836 20292 3845
rect 19972 3834 19996 3836
rect 20052 3834 20076 3836
rect 20132 3834 20156 3836
rect 20212 3834 20236 3836
rect 19972 3782 19982 3834
rect 20226 3782 20236 3834
rect 19972 3780 19996 3782
rect 20052 3780 20076 3782
rect 20132 3780 20156 3782
rect 20212 3780 20236 3782
rect 19916 3771 20292 3780
rect 20656 3292 21032 3301
rect 20712 3290 20736 3292
rect 20792 3290 20816 3292
rect 20872 3290 20896 3292
rect 20952 3290 20976 3292
rect 20712 3238 20722 3290
rect 20966 3238 20976 3290
rect 20712 3236 20736 3238
rect 20792 3236 20816 3238
rect 20872 3236 20896 3238
rect 20952 3236 20976 3238
rect 20656 3227 21032 3236
rect 18064 2746 18276 2774
rect 18248 2446 18276 2746
rect 19916 2748 20292 2757
rect 19972 2746 19996 2748
rect 20052 2746 20076 2748
rect 20132 2746 20156 2748
rect 20212 2746 20236 2748
rect 19972 2694 19982 2746
rect 20226 2694 20236 2746
rect 19972 2692 19996 2694
rect 20052 2692 20076 2694
rect 20132 2692 20156 2694
rect 20212 2692 20236 2694
rect 19916 2683 20292 2692
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 17040 2440 17092 2446
rect 17040 2382 17092 2388
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 12164 2372 12216 2378
rect 12164 2314 12216 2320
rect 12900 2372 12952 2378
rect 12900 2314 12952 2320
rect 13544 2372 13596 2378
rect 13544 2314 13596 2320
rect 17316 2372 17368 2378
rect 17316 2314 17368 2320
rect 18052 2372 18104 2378
rect 18052 2314 18104 2320
rect 12176 1170 12204 2314
rect 12176 1142 12296 1170
rect 12268 800 12296 1142
rect 12912 800 12940 2314
rect 13556 800 13584 2314
rect 14656 2204 15032 2213
rect 14712 2202 14736 2204
rect 14792 2202 14816 2204
rect 14872 2202 14896 2204
rect 14952 2202 14976 2204
rect 14712 2150 14722 2202
rect 14966 2150 14976 2202
rect 14712 2148 14736 2150
rect 14792 2148 14816 2150
rect 14872 2148 14896 2150
rect 14952 2148 14976 2150
rect 14656 2139 15032 2148
rect 17328 1170 17356 2314
rect 17328 1142 17448 1170
rect 17420 800 17448 1142
rect 18064 800 18092 2314
rect 20656 2204 21032 2213
rect 20712 2202 20736 2204
rect 20792 2202 20816 2204
rect 20872 2202 20896 2204
rect 20952 2202 20976 2204
rect 20712 2150 20722 2202
rect 20966 2150 20976 2202
rect 20712 2148 20736 2150
rect 20792 2148 20816 2150
rect 20872 2148 20896 2150
rect 20952 2148 20976 2150
rect 20656 2139 21032 2148
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 17406 0 17462 800
rect 18050 0 18106 800
<< via2 >>
rect 1916 24506 1972 24508
rect 1996 24506 2052 24508
rect 2076 24506 2132 24508
rect 2156 24506 2212 24508
rect 2236 24506 2292 24508
rect 1916 24454 1918 24506
rect 1918 24454 1970 24506
rect 1970 24454 1972 24506
rect 1996 24454 2034 24506
rect 2034 24454 2046 24506
rect 2046 24454 2052 24506
rect 2076 24454 2098 24506
rect 2098 24454 2110 24506
rect 2110 24454 2132 24506
rect 2156 24454 2162 24506
rect 2162 24454 2174 24506
rect 2174 24454 2212 24506
rect 2236 24454 2238 24506
rect 2238 24454 2290 24506
rect 2290 24454 2292 24506
rect 1916 24452 1972 24454
rect 1996 24452 2052 24454
rect 2076 24452 2132 24454
rect 2156 24452 2212 24454
rect 2236 24452 2292 24454
rect 7916 24506 7972 24508
rect 7996 24506 8052 24508
rect 8076 24506 8132 24508
rect 8156 24506 8212 24508
rect 8236 24506 8292 24508
rect 7916 24454 7918 24506
rect 7918 24454 7970 24506
rect 7970 24454 7972 24506
rect 7996 24454 8034 24506
rect 8034 24454 8046 24506
rect 8046 24454 8052 24506
rect 8076 24454 8098 24506
rect 8098 24454 8110 24506
rect 8110 24454 8132 24506
rect 8156 24454 8162 24506
rect 8162 24454 8174 24506
rect 8174 24454 8212 24506
rect 8236 24454 8238 24506
rect 8238 24454 8290 24506
rect 8290 24454 8292 24506
rect 7916 24452 7972 24454
rect 7996 24452 8052 24454
rect 8076 24452 8132 24454
rect 8156 24452 8212 24454
rect 8236 24452 8292 24454
rect 13916 24506 13972 24508
rect 13996 24506 14052 24508
rect 14076 24506 14132 24508
rect 14156 24506 14212 24508
rect 14236 24506 14292 24508
rect 13916 24454 13918 24506
rect 13918 24454 13970 24506
rect 13970 24454 13972 24506
rect 13996 24454 14034 24506
rect 14034 24454 14046 24506
rect 14046 24454 14052 24506
rect 14076 24454 14098 24506
rect 14098 24454 14110 24506
rect 14110 24454 14132 24506
rect 14156 24454 14162 24506
rect 14162 24454 14174 24506
rect 14174 24454 14212 24506
rect 14236 24454 14238 24506
rect 14238 24454 14290 24506
rect 14290 24454 14292 24506
rect 13916 24452 13972 24454
rect 13996 24452 14052 24454
rect 14076 24452 14132 24454
rect 14156 24452 14212 24454
rect 14236 24452 14292 24454
rect 19916 24506 19972 24508
rect 19996 24506 20052 24508
rect 20076 24506 20132 24508
rect 20156 24506 20212 24508
rect 20236 24506 20292 24508
rect 19916 24454 19918 24506
rect 19918 24454 19970 24506
rect 19970 24454 19972 24506
rect 19996 24454 20034 24506
rect 20034 24454 20046 24506
rect 20046 24454 20052 24506
rect 20076 24454 20098 24506
rect 20098 24454 20110 24506
rect 20110 24454 20132 24506
rect 20156 24454 20162 24506
rect 20162 24454 20174 24506
rect 20174 24454 20212 24506
rect 20236 24454 20238 24506
rect 20238 24454 20290 24506
rect 20290 24454 20292 24506
rect 19916 24452 19972 24454
rect 19996 24452 20052 24454
rect 20076 24452 20132 24454
rect 20156 24452 20212 24454
rect 20236 24452 20292 24454
rect 2656 23962 2712 23964
rect 2736 23962 2792 23964
rect 2816 23962 2872 23964
rect 2896 23962 2952 23964
rect 2976 23962 3032 23964
rect 2656 23910 2658 23962
rect 2658 23910 2710 23962
rect 2710 23910 2712 23962
rect 2736 23910 2774 23962
rect 2774 23910 2786 23962
rect 2786 23910 2792 23962
rect 2816 23910 2838 23962
rect 2838 23910 2850 23962
rect 2850 23910 2872 23962
rect 2896 23910 2902 23962
rect 2902 23910 2914 23962
rect 2914 23910 2952 23962
rect 2976 23910 2978 23962
rect 2978 23910 3030 23962
rect 3030 23910 3032 23962
rect 2656 23908 2712 23910
rect 2736 23908 2792 23910
rect 2816 23908 2872 23910
rect 2896 23908 2952 23910
rect 2976 23908 3032 23910
rect 1916 23418 1972 23420
rect 1996 23418 2052 23420
rect 2076 23418 2132 23420
rect 2156 23418 2212 23420
rect 2236 23418 2292 23420
rect 1916 23366 1918 23418
rect 1918 23366 1970 23418
rect 1970 23366 1972 23418
rect 1996 23366 2034 23418
rect 2034 23366 2046 23418
rect 2046 23366 2052 23418
rect 2076 23366 2098 23418
rect 2098 23366 2110 23418
rect 2110 23366 2132 23418
rect 2156 23366 2162 23418
rect 2162 23366 2174 23418
rect 2174 23366 2212 23418
rect 2236 23366 2238 23418
rect 2238 23366 2290 23418
rect 2290 23366 2292 23418
rect 1916 23364 1972 23366
rect 1996 23364 2052 23366
rect 2076 23364 2132 23366
rect 2156 23364 2212 23366
rect 2236 23364 2292 23366
rect 2656 22874 2712 22876
rect 2736 22874 2792 22876
rect 2816 22874 2872 22876
rect 2896 22874 2952 22876
rect 2976 22874 3032 22876
rect 2656 22822 2658 22874
rect 2658 22822 2710 22874
rect 2710 22822 2712 22874
rect 2736 22822 2774 22874
rect 2774 22822 2786 22874
rect 2786 22822 2792 22874
rect 2816 22822 2838 22874
rect 2838 22822 2850 22874
rect 2850 22822 2872 22874
rect 2896 22822 2902 22874
rect 2902 22822 2914 22874
rect 2914 22822 2952 22874
rect 2976 22822 2978 22874
rect 2978 22822 3030 22874
rect 3030 22822 3032 22874
rect 2656 22820 2712 22822
rect 2736 22820 2792 22822
rect 2816 22820 2872 22822
rect 2896 22820 2952 22822
rect 2976 22820 3032 22822
rect 1916 22330 1972 22332
rect 1996 22330 2052 22332
rect 2076 22330 2132 22332
rect 2156 22330 2212 22332
rect 2236 22330 2292 22332
rect 1916 22278 1918 22330
rect 1918 22278 1970 22330
rect 1970 22278 1972 22330
rect 1996 22278 2034 22330
rect 2034 22278 2046 22330
rect 2046 22278 2052 22330
rect 2076 22278 2098 22330
rect 2098 22278 2110 22330
rect 2110 22278 2132 22330
rect 2156 22278 2162 22330
rect 2162 22278 2174 22330
rect 2174 22278 2212 22330
rect 2236 22278 2238 22330
rect 2238 22278 2290 22330
rect 2290 22278 2292 22330
rect 1916 22276 1972 22278
rect 1996 22276 2052 22278
rect 2076 22276 2132 22278
rect 2156 22276 2212 22278
rect 2236 22276 2292 22278
rect 2656 21786 2712 21788
rect 2736 21786 2792 21788
rect 2816 21786 2872 21788
rect 2896 21786 2952 21788
rect 2976 21786 3032 21788
rect 2656 21734 2658 21786
rect 2658 21734 2710 21786
rect 2710 21734 2712 21786
rect 2736 21734 2774 21786
rect 2774 21734 2786 21786
rect 2786 21734 2792 21786
rect 2816 21734 2838 21786
rect 2838 21734 2850 21786
rect 2850 21734 2872 21786
rect 2896 21734 2902 21786
rect 2902 21734 2914 21786
rect 2914 21734 2952 21786
rect 2976 21734 2978 21786
rect 2978 21734 3030 21786
rect 3030 21734 3032 21786
rect 2656 21732 2712 21734
rect 2736 21732 2792 21734
rect 2816 21732 2872 21734
rect 2896 21732 2952 21734
rect 2976 21732 3032 21734
rect 1916 21242 1972 21244
rect 1996 21242 2052 21244
rect 2076 21242 2132 21244
rect 2156 21242 2212 21244
rect 2236 21242 2292 21244
rect 1916 21190 1918 21242
rect 1918 21190 1970 21242
rect 1970 21190 1972 21242
rect 1996 21190 2034 21242
rect 2034 21190 2046 21242
rect 2046 21190 2052 21242
rect 2076 21190 2098 21242
rect 2098 21190 2110 21242
rect 2110 21190 2132 21242
rect 2156 21190 2162 21242
rect 2162 21190 2174 21242
rect 2174 21190 2212 21242
rect 2236 21190 2238 21242
rect 2238 21190 2290 21242
rect 2290 21190 2292 21242
rect 1916 21188 1972 21190
rect 1996 21188 2052 21190
rect 2076 21188 2132 21190
rect 2156 21188 2212 21190
rect 2236 21188 2292 21190
rect 2656 20698 2712 20700
rect 2736 20698 2792 20700
rect 2816 20698 2872 20700
rect 2896 20698 2952 20700
rect 2976 20698 3032 20700
rect 2656 20646 2658 20698
rect 2658 20646 2710 20698
rect 2710 20646 2712 20698
rect 2736 20646 2774 20698
rect 2774 20646 2786 20698
rect 2786 20646 2792 20698
rect 2816 20646 2838 20698
rect 2838 20646 2850 20698
rect 2850 20646 2872 20698
rect 2896 20646 2902 20698
rect 2902 20646 2914 20698
rect 2914 20646 2952 20698
rect 2976 20646 2978 20698
rect 2978 20646 3030 20698
rect 3030 20646 3032 20698
rect 2656 20644 2712 20646
rect 2736 20644 2792 20646
rect 2816 20644 2872 20646
rect 2896 20644 2952 20646
rect 2976 20644 3032 20646
rect 1916 20154 1972 20156
rect 1996 20154 2052 20156
rect 2076 20154 2132 20156
rect 2156 20154 2212 20156
rect 2236 20154 2292 20156
rect 1916 20102 1918 20154
rect 1918 20102 1970 20154
rect 1970 20102 1972 20154
rect 1996 20102 2034 20154
rect 2034 20102 2046 20154
rect 2046 20102 2052 20154
rect 2076 20102 2098 20154
rect 2098 20102 2110 20154
rect 2110 20102 2132 20154
rect 2156 20102 2162 20154
rect 2162 20102 2174 20154
rect 2174 20102 2212 20154
rect 2236 20102 2238 20154
rect 2238 20102 2290 20154
rect 2290 20102 2292 20154
rect 1916 20100 1972 20102
rect 1996 20100 2052 20102
rect 2076 20100 2132 20102
rect 2156 20100 2212 20102
rect 2236 20100 2292 20102
rect 3790 19760 3846 19816
rect 2656 19610 2712 19612
rect 2736 19610 2792 19612
rect 2816 19610 2872 19612
rect 2896 19610 2952 19612
rect 2976 19610 3032 19612
rect 2656 19558 2658 19610
rect 2658 19558 2710 19610
rect 2710 19558 2712 19610
rect 2736 19558 2774 19610
rect 2774 19558 2786 19610
rect 2786 19558 2792 19610
rect 2816 19558 2838 19610
rect 2838 19558 2850 19610
rect 2850 19558 2872 19610
rect 2896 19558 2902 19610
rect 2902 19558 2914 19610
rect 2914 19558 2952 19610
rect 2976 19558 2978 19610
rect 2978 19558 3030 19610
rect 3030 19558 3032 19610
rect 2656 19556 2712 19558
rect 2736 19556 2792 19558
rect 2816 19556 2872 19558
rect 2896 19556 2952 19558
rect 2976 19556 3032 19558
rect 1916 19066 1972 19068
rect 1996 19066 2052 19068
rect 2076 19066 2132 19068
rect 2156 19066 2212 19068
rect 2236 19066 2292 19068
rect 1916 19014 1918 19066
rect 1918 19014 1970 19066
rect 1970 19014 1972 19066
rect 1996 19014 2034 19066
rect 2034 19014 2046 19066
rect 2046 19014 2052 19066
rect 2076 19014 2098 19066
rect 2098 19014 2110 19066
rect 2110 19014 2132 19066
rect 2156 19014 2162 19066
rect 2162 19014 2174 19066
rect 2174 19014 2212 19066
rect 2236 19014 2238 19066
rect 2238 19014 2290 19066
rect 2290 19014 2292 19066
rect 1916 19012 1972 19014
rect 1996 19012 2052 19014
rect 2076 19012 2132 19014
rect 2156 19012 2212 19014
rect 2236 19012 2292 19014
rect 2656 18522 2712 18524
rect 2736 18522 2792 18524
rect 2816 18522 2872 18524
rect 2896 18522 2952 18524
rect 2976 18522 3032 18524
rect 2656 18470 2658 18522
rect 2658 18470 2710 18522
rect 2710 18470 2712 18522
rect 2736 18470 2774 18522
rect 2774 18470 2786 18522
rect 2786 18470 2792 18522
rect 2816 18470 2838 18522
rect 2838 18470 2850 18522
rect 2850 18470 2872 18522
rect 2896 18470 2902 18522
rect 2902 18470 2914 18522
rect 2914 18470 2952 18522
rect 2976 18470 2978 18522
rect 2978 18470 3030 18522
rect 3030 18470 3032 18522
rect 2656 18468 2712 18470
rect 2736 18468 2792 18470
rect 2816 18468 2872 18470
rect 2896 18468 2952 18470
rect 2976 18468 3032 18470
rect 1916 17978 1972 17980
rect 1996 17978 2052 17980
rect 2076 17978 2132 17980
rect 2156 17978 2212 17980
rect 2236 17978 2292 17980
rect 1916 17926 1918 17978
rect 1918 17926 1970 17978
rect 1970 17926 1972 17978
rect 1996 17926 2034 17978
rect 2034 17926 2046 17978
rect 2046 17926 2052 17978
rect 2076 17926 2098 17978
rect 2098 17926 2110 17978
rect 2110 17926 2132 17978
rect 2156 17926 2162 17978
rect 2162 17926 2174 17978
rect 2174 17926 2212 17978
rect 2236 17926 2238 17978
rect 2238 17926 2290 17978
rect 2290 17926 2292 17978
rect 1916 17924 1972 17926
rect 1996 17924 2052 17926
rect 2076 17924 2132 17926
rect 2156 17924 2212 17926
rect 2236 17924 2292 17926
rect 2656 17434 2712 17436
rect 2736 17434 2792 17436
rect 2816 17434 2872 17436
rect 2896 17434 2952 17436
rect 2976 17434 3032 17436
rect 2656 17382 2658 17434
rect 2658 17382 2710 17434
rect 2710 17382 2712 17434
rect 2736 17382 2774 17434
rect 2774 17382 2786 17434
rect 2786 17382 2792 17434
rect 2816 17382 2838 17434
rect 2838 17382 2850 17434
rect 2850 17382 2872 17434
rect 2896 17382 2902 17434
rect 2902 17382 2914 17434
rect 2914 17382 2952 17434
rect 2976 17382 2978 17434
rect 2978 17382 3030 17434
rect 3030 17382 3032 17434
rect 2656 17380 2712 17382
rect 2736 17380 2792 17382
rect 2816 17380 2872 17382
rect 2896 17380 2952 17382
rect 2976 17380 3032 17382
rect 938 17076 940 17096
rect 940 17076 992 17096
rect 992 17076 994 17096
rect 938 17040 994 17076
rect 1916 16890 1972 16892
rect 1996 16890 2052 16892
rect 2076 16890 2132 16892
rect 2156 16890 2212 16892
rect 2236 16890 2292 16892
rect 1916 16838 1918 16890
rect 1918 16838 1970 16890
rect 1970 16838 1972 16890
rect 1996 16838 2034 16890
rect 2034 16838 2046 16890
rect 2046 16838 2052 16890
rect 2076 16838 2098 16890
rect 2098 16838 2110 16890
rect 2110 16838 2132 16890
rect 2156 16838 2162 16890
rect 2162 16838 2174 16890
rect 2174 16838 2212 16890
rect 2236 16838 2238 16890
rect 2238 16838 2290 16890
rect 2290 16838 2292 16890
rect 1916 16836 1972 16838
rect 1996 16836 2052 16838
rect 2076 16836 2132 16838
rect 2156 16836 2212 16838
rect 2236 16836 2292 16838
rect 938 15680 994 15736
rect 938 13640 994 13696
rect 938 12280 994 12336
rect 1858 15952 1914 16008
rect 1916 15802 1972 15804
rect 1996 15802 2052 15804
rect 2076 15802 2132 15804
rect 2156 15802 2212 15804
rect 2236 15802 2292 15804
rect 1916 15750 1918 15802
rect 1918 15750 1970 15802
rect 1970 15750 1972 15802
rect 1996 15750 2034 15802
rect 2034 15750 2046 15802
rect 2046 15750 2052 15802
rect 2076 15750 2098 15802
rect 2098 15750 2110 15802
rect 2110 15750 2132 15802
rect 2156 15750 2162 15802
rect 2162 15750 2174 15802
rect 2174 15750 2212 15802
rect 2236 15750 2238 15802
rect 2238 15750 2290 15802
rect 2290 15750 2292 15802
rect 1916 15748 1972 15750
rect 1996 15748 2052 15750
rect 2076 15748 2132 15750
rect 2156 15748 2212 15750
rect 2236 15748 2292 15750
rect 2226 15544 2282 15600
rect 1306 13096 1362 13152
rect 1214 7928 1270 7984
rect 1916 14714 1972 14716
rect 1996 14714 2052 14716
rect 2076 14714 2132 14716
rect 2156 14714 2212 14716
rect 2236 14714 2292 14716
rect 1916 14662 1918 14714
rect 1918 14662 1970 14714
rect 1970 14662 1972 14714
rect 1996 14662 2034 14714
rect 2034 14662 2046 14714
rect 2046 14662 2052 14714
rect 2076 14662 2098 14714
rect 2098 14662 2110 14714
rect 2110 14662 2132 14714
rect 2156 14662 2162 14714
rect 2162 14662 2174 14714
rect 2174 14662 2212 14714
rect 2236 14662 2238 14714
rect 2238 14662 2290 14714
rect 2290 14662 2292 14714
rect 1916 14660 1972 14662
rect 1996 14660 2052 14662
rect 2076 14660 2132 14662
rect 2156 14660 2212 14662
rect 2236 14660 2292 14662
rect 1916 13626 1972 13628
rect 1996 13626 2052 13628
rect 2076 13626 2132 13628
rect 2156 13626 2212 13628
rect 2236 13626 2292 13628
rect 1916 13574 1918 13626
rect 1918 13574 1970 13626
rect 1970 13574 1972 13626
rect 1996 13574 2034 13626
rect 2034 13574 2046 13626
rect 2046 13574 2052 13626
rect 2076 13574 2098 13626
rect 2098 13574 2110 13626
rect 2110 13574 2132 13626
rect 2156 13574 2162 13626
rect 2162 13574 2174 13626
rect 2174 13574 2212 13626
rect 2236 13574 2238 13626
rect 2238 13574 2290 13626
rect 2290 13574 2292 13626
rect 1916 13572 1972 13574
rect 1996 13572 2052 13574
rect 2076 13572 2132 13574
rect 2156 13572 2212 13574
rect 2236 13572 2292 13574
rect 1916 12538 1972 12540
rect 1996 12538 2052 12540
rect 2076 12538 2132 12540
rect 2156 12538 2212 12540
rect 2236 12538 2292 12540
rect 1916 12486 1918 12538
rect 1918 12486 1970 12538
rect 1970 12486 1972 12538
rect 1996 12486 2034 12538
rect 2034 12486 2046 12538
rect 2046 12486 2052 12538
rect 2076 12486 2098 12538
rect 2098 12486 2110 12538
rect 2110 12486 2132 12538
rect 2156 12486 2162 12538
rect 2162 12486 2174 12538
rect 2174 12486 2212 12538
rect 2236 12486 2238 12538
rect 2238 12486 2290 12538
rect 2290 12486 2292 12538
rect 1916 12484 1972 12486
rect 1996 12484 2052 12486
rect 2076 12484 2132 12486
rect 2156 12484 2212 12486
rect 2236 12484 2292 12486
rect 1766 11620 1822 11656
rect 1766 11600 1768 11620
rect 1768 11600 1820 11620
rect 1820 11600 1822 11620
rect 1916 11450 1972 11452
rect 1996 11450 2052 11452
rect 2076 11450 2132 11452
rect 2156 11450 2212 11452
rect 2236 11450 2292 11452
rect 1916 11398 1918 11450
rect 1918 11398 1970 11450
rect 1970 11398 1972 11450
rect 1996 11398 2034 11450
rect 2034 11398 2046 11450
rect 2046 11398 2052 11450
rect 2076 11398 2098 11450
rect 2098 11398 2110 11450
rect 2110 11398 2132 11450
rect 2156 11398 2162 11450
rect 2162 11398 2174 11450
rect 2174 11398 2212 11450
rect 2236 11398 2238 11450
rect 2238 11398 2290 11450
rect 2290 11398 2292 11450
rect 1916 11396 1972 11398
rect 1996 11396 2052 11398
rect 2076 11396 2132 11398
rect 2156 11396 2212 11398
rect 2236 11396 2292 11398
rect 2656 16346 2712 16348
rect 2736 16346 2792 16348
rect 2816 16346 2872 16348
rect 2896 16346 2952 16348
rect 2976 16346 3032 16348
rect 2656 16294 2658 16346
rect 2658 16294 2710 16346
rect 2710 16294 2712 16346
rect 2736 16294 2774 16346
rect 2774 16294 2786 16346
rect 2786 16294 2792 16346
rect 2816 16294 2838 16346
rect 2838 16294 2850 16346
rect 2850 16294 2872 16346
rect 2896 16294 2902 16346
rect 2902 16294 2914 16346
rect 2914 16294 2952 16346
rect 2976 16294 2978 16346
rect 2978 16294 3030 16346
rect 3030 16294 3032 16346
rect 2656 16292 2712 16294
rect 2736 16292 2792 16294
rect 2816 16292 2872 16294
rect 2896 16292 2952 16294
rect 2976 16292 3032 16294
rect 1674 7792 1730 7848
rect 1916 10362 1972 10364
rect 1996 10362 2052 10364
rect 2076 10362 2132 10364
rect 2156 10362 2212 10364
rect 2236 10362 2292 10364
rect 1916 10310 1918 10362
rect 1918 10310 1970 10362
rect 1970 10310 1972 10362
rect 1996 10310 2034 10362
rect 2034 10310 2046 10362
rect 2046 10310 2052 10362
rect 2076 10310 2098 10362
rect 2098 10310 2110 10362
rect 2110 10310 2132 10362
rect 2156 10310 2162 10362
rect 2162 10310 2174 10362
rect 2174 10310 2212 10362
rect 2236 10310 2238 10362
rect 2238 10310 2290 10362
rect 2290 10310 2292 10362
rect 1916 10308 1972 10310
rect 1996 10308 2052 10310
rect 2076 10308 2132 10310
rect 2156 10308 2212 10310
rect 2236 10308 2292 10310
rect 2226 9580 2282 9616
rect 2226 9560 2228 9580
rect 2228 9560 2280 9580
rect 2280 9560 2282 9580
rect 1916 9274 1972 9276
rect 1996 9274 2052 9276
rect 2076 9274 2132 9276
rect 2156 9274 2212 9276
rect 2236 9274 2292 9276
rect 1916 9222 1918 9274
rect 1918 9222 1970 9274
rect 1970 9222 1972 9274
rect 1996 9222 2034 9274
rect 2034 9222 2046 9274
rect 2046 9222 2052 9274
rect 2076 9222 2098 9274
rect 2098 9222 2110 9274
rect 2110 9222 2132 9274
rect 2156 9222 2162 9274
rect 2162 9222 2174 9274
rect 2174 9222 2212 9274
rect 2236 9222 2238 9274
rect 2238 9222 2290 9274
rect 2290 9222 2292 9274
rect 1916 9220 1972 9222
rect 1996 9220 2052 9222
rect 2076 9220 2132 9222
rect 2156 9220 2212 9222
rect 2236 9220 2292 9222
rect 2594 15408 2650 15464
rect 2656 15258 2712 15260
rect 2736 15258 2792 15260
rect 2816 15258 2872 15260
rect 2896 15258 2952 15260
rect 2976 15258 3032 15260
rect 2656 15206 2658 15258
rect 2658 15206 2710 15258
rect 2710 15206 2712 15258
rect 2736 15206 2774 15258
rect 2774 15206 2786 15258
rect 2786 15206 2792 15258
rect 2816 15206 2838 15258
rect 2838 15206 2850 15258
rect 2850 15206 2872 15258
rect 2896 15206 2902 15258
rect 2902 15206 2914 15258
rect 2914 15206 2952 15258
rect 2976 15206 2978 15258
rect 2978 15206 3030 15258
rect 3030 15206 3032 15258
rect 2656 15204 2712 15206
rect 2736 15204 2792 15206
rect 2816 15204 2872 15206
rect 2896 15204 2952 15206
rect 2976 15204 3032 15206
rect 3422 17040 3478 17096
rect 3606 16088 3662 16144
rect 3606 15544 3662 15600
rect 2656 14170 2712 14172
rect 2736 14170 2792 14172
rect 2816 14170 2872 14172
rect 2896 14170 2952 14172
rect 2976 14170 3032 14172
rect 2656 14118 2658 14170
rect 2658 14118 2710 14170
rect 2710 14118 2712 14170
rect 2736 14118 2774 14170
rect 2774 14118 2786 14170
rect 2786 14118 2792 14170
rect 2816 14118 2838 14170
rect 2838 14118 2850 14170
rect 2850 14118 2872 14170
rect 2896 14118 2902 14170
rect 2902 14118 2914 14170
rect 2914 14118 2952 14170
rect 2976 14118 2978 14170
rect 2978 14118 3030 14170
rect 3030 14118 3032 14170
rect 2656 14116 2712 14118
rect 2736 14116 2792 14118
rect 2816 14116 2872 14118
rect 2896 14116 2952 14118
rect 2976 14116 3032 14118
rect 3882 16632 3938 16688
rect 3790 13368 3846 13424
rect 4250 15408 4306 15464
rect 2656 13082 2712 13084
rect 2736 13082 2792 13084
rect 2816 13082 2872 13084
rect 2896 13082 2952 13084
rect 2976 13082 3032 13084
rect 2656 13030 2658 13082
rect 2658 13030 2710 13082
rect 2710 13030 2712 13082
rect 2736 13030 2774 13082
rect 2774 13030 2786 13082
rect 2786 13030 2792 13082
rect 2816 13030 2838 13082
rect 2838 13030 2850 13082
rect 2850 13030 2872 13082
rect 2896 13030 2902 13082
rect 2902 13030 2914 13082
rect 2914 13030 2952 13082
rect 2976 13030 2978 13082
rect 2978 13030 3030 13082
rect 3030 13030 3032 13082
rect 2656 13028 2712 13030
rect 2736 13028 2792 13030
rect 2816 13028 2872 13030
rect 2896 13028 2952 13030
rect 2976 13028 3032 13030
rect 2656 11994 2712 11996
rect 2736 11994 2792 11996
rect 2816 11994 2872 11996
rect 2896 11994 2952 11996
rect 2976 11994 3032 11996
rect 2656 11942 2658 11994
rect 2658 11942 2710 11994
rect 2710 11942 2712 11994
rect 2736 11942 2774 11994
rect 2774 11942 2786 11994
rect 2786 11942 2792 11994
rect 2816 11942 2838 11994
rect 2838 11942 2850 11994
rect 2850 11942 2872 11994
rect 2896 11942 2902 11994
rect 2902 11942 2914 11994
rect 2914 11942 2952 11994
rect 2976 11942 2978 11994
rect 2978 11942 3030 11994
rect 3030 11942 3032 11994
rect 2656 11940 2712 11942
rect 2736 11940 2792 11942
rect 2816 11940 2872 11942
rect 2896 11940 2952 11942
rect 2976 11940 3032 11942
rect 2656 10906 2712 10908
rect 2736 10906 2792 10908
rect 2816 10906 2872 10908
rect 2896 10906 2952 10908
rect 2976 10906 3032 10908
rect 2656 10854 2658 10906
rect 2658 10854 2710 10906
rect 2710 10854 2712 10906
rect 2736 10854 2774 10906
rect 2774 10854 2786 10906
rect 2786 10854 2792 10906
rect 2816 10854 2838 10906
rect 2838 10854 2850 10906
rect 2850 10854 2872 10906
rect 2896 10854 2902 10906
rect 2902 10854 2914 10906
rect 2914 10854 2952 10906
rect 2976 10854 2978 10906
rect 2978 10854 3030 10906
rect 3030 10854 3032 10906
rect 2656 10852 2712 10854
rect 2736 10852 2792 10854
rect 2816 10852 2872 10854
rect 2896 10852 2952 10854
rect 2976 10852 3032 10854
rect 2656 9818 2712 9820
rect 2736 9818 2792 9820
rect 2816 9818 2872 9820
rect 2896 9818 2952 9820
rect 2976 9818 3032 9820
rect 2656 9766 2658 9818
rect 2658 9766 2710 9818
rect 2710 9766 2712 9818
rect 2736 9766 2774 9818
rect 2774 9766 2786 9818
rect 2786 9766 2792 9818
rect 2816 9766 2838 9818
rect 2838 9766 2850 9818
rect 2850 9766 2872 9818
rect 2896 9766 2902 9818
rect 2902 9766 2914 9818
rect 2914 9766 2952 9818
rect 2976 9766 2978 9818
rect 2978 9766 3030 9818
rect 3030 9766 3032 9818
rect 2656 9764 2712 9766
rect 2736 9764 2792 9766
rect 2816 9764 2872 9766
rect 2896 9764 2952 9766
rect 2976 9764 3032 9766
rect 2410 9444 2466 9480
rect 2410 9424 2412 9444
rect 2412 9424 2464 9444
rect 2464 9424 2466 9444
rect 2656 8730 2712 8732
rect 2736 8730 2792 8732
rect 2816 8730 2872 8732
rect 2896 8730 2952 8732
rect 2976 8730 3032 8732
rect 2656 8678 2658 8730
rect 2658 8678 2710 8730
rect 2710 8678 2712 8730
rect 2736 8678 2774 8730
rect 2774 8678 2786 8730
rect 2786 8678 2792 8730
rect 2816 8678 2838 8730
rect 2838 8678 2850 8730
rect 2850 8678 2872 8730
rect 2896 8678 2902 8730
rect 2902 8678 2914 8730
rect 2914 8678 2952 8730
rect 2976 8678 2978 8730
rect 2978 8678 3030 8730
rect 3030 8678 3032 8730
rect 2656 8676 2712 8678
rect 2736 8676 2792 8678
rect 2816 8676 2872 8678
rect 2896 8676 2952 8678
rect 2976 8676 3032 8678
rect 1916 8186 1972 8188
rect 1996 8186 2052 8188
rect 2076 8186 2132 8188
rect 2156 8186 2212 8188
rect 2236 8186 2292 8188
rect 1916 8134 1918 8186
rect 1918 8134 1970 8186
rect 1970 8134 1972 8186
rect 1996 8134 2034 8186
rect 2034 8134 2046 8186
rect 2046 8134 2052 8186
rect 2076 8134 2098 8186
rect 2098 8134 2110 8186
rect 2110 8134 2132 8186
rect 2156 8134 2162 8186
rect 2162 8134 2174 8186
rect 2174 8134 2212 8186
rect 2236 8134 2238 8186
rect 2238 8134 2290 8186
rect 2290 8134 2292 8186
rect 1916 8132 1972 8134
rect 1996 8132 2052 8134
rect 2076 8132 2132 8134
rect 2156 8132 2212 8134
rect 2236 8132 2292 8134
rect 1916 7098 1972 7100
rect 1996 7098 2052 7100
rect 2076 7098 2132 7100
rect 2156 7098 2212 7100
rect 2236 7098 2292 7100
rect 1916 7046 1918 7098
rect 1918 7046 1970 7098
rect 1970 7046 1972 7098
rect 1996 7046 2034 7098
rect 2034 7046 2046 7098
rect 2046 7046 2052 7098
rect 2076 7046 2098 7098
rect 2098 7046 2110 7098
rect 2110 7046 2132 7098
rect 2156 7046 2162 7098
rect 2162 7046 2174 7098
rect 2174 7046 2212 7098
rect 2236 7046 2238 7098
rect 2238 7046 2290 7098
rect 2290 7046 2292 7098
rect 1916 7044 1972 7046
rect 1996 7044 2052 7046
rect 2076 7044 2132 7046
rect 2156 7044 2212 7046
rect 2236 7044 2292 7046
rect 1916 6010 1972 6012
rect 1996 6010 2052 6012
rect 2076 6010 2132 6012
rect 2156 6010 2212 6012
rect 2236 6010 2292 6012
rect 1916 5958 1918 6010
rect 1918 5958 1970 6010
rect 1970 5958 1972 6010
rect 1996 5958 2034 6010
rect 2034 5958 2046 6010
rect 2046 5958 2052 6010
rect 2076 5958 2098 6010
rect 2098 5958 2110 6010
rect 2110 5958 2132 6010
rect 2156 5958 2162 6010
rect 2162 5958 2174 6010
rect 2174 5958 2212 6010
rect 2236 5958 2238 6010
rect 2238 5958 2290 6010
rect 2290 5958 2292 6010
rect 1916 5956 1972 5958
rect 1996 5956 2052 5958
rect 2076 5956 2132 5958
rect 2156 5956 2212 5958
rect 2236 5956 2292 5958
rect 2226 5752 2282 5808
rect 2594 7928 2650 7984
rect 2656 7642 2712 7644
rect 2736 7642 2792 7644
rect 2816 7642 2872 7644
rect 2896 7642 2952 7644
rect 2976 7642 3032 7644
rect 2656 7590 2658 7642
rect 2658 7590 2710 7642
rect 2710 7590 2712 7642
rect 2736 7590 2774 7642
rect 2774 7590 2786 7642
rect 2786 7590 2792 7642
rect 2816 7590 2838 7642
rect 2838 7590 2850 7642
rect 2850 7590 2872 7642
rect 2896 7590 2902 7642
rect 2902 7590 2914 7642
rect 2914 7590 2952 7642
rect 2976 7590 2978 7642
rect 2978 7590 3030 7642
rect 3030 7590 3032 7642
rect 2656 7588 2712 7590
rect 2736 7588 2792 7590
rect 2816 7588 2872 7590
rect 2896 7588 2952 7590
rect 2976 7588 3032 7590
rect 3790 12824 3846 12880
rect 3054 7284 3056 7304
rect 3056 7284 3108 7304
rect 3108 7284 3110 7304
rect 3054 7248 3110 7284
rect 2686 7112 2742 7168
rect 2410 6024 2466 6080
rect 2778 6976 2834 7032
rect 3054 6876 3056 6896
rect 3056 6876 3108 6896
rect 3108 6876 3110 6896
rect 3054 6840 3110 6876
rect 2656 6554 2712 6556
rect 2736 6554 2792 6556
rect 2816 6554 2872 6556
rect 2896 6554 2952 6556
rect 2976 6554 3032 6556
rect 2656 6502 2658 6554
rect 2658 6502 2710 6554
rect 2710 6502 2712 6554
rect 2736 6502 2774 6554
rect 2774 6502 2786 6554
rect 2786 6502 2792 6554
rect 2816 6502 2838 6554
rect 2838 6502 2850 6554
rect 2850 6502 2872 6554
rect 2896 6502 2902 6554
rect 2902 6502 2914 6554
rect 2914 6502 2952 6554
rect 2976 6502 2978 6554
rect 2978 6502 3030 6554
rect 3030 6502 3032 6554
rect 2656 6500 2712 6502
rect 2736 6500 2792 6502
rect 2816 6500 2872 6502
rect 2896 6500 2952 6502
rect 2976 6500 3032 6502
rect 3054 6296 3110 6352
rect 3054 6196 3056 6216
rect 3056 6196 3108 6216
rect 3108 6196 3110 6216
rect 3054 6160 3110 6196
rect 3054 5888 3110 5944
rect 2870 5616 2926 5672
rect 2656 5466 2712 5468
rect 2736 5466 2792 5468
rect 2816 5466 2872 5468
rect 2896 5466 2952 5468
rect 2976 5466 3032 5468
rect 2656 5414 2658 5466
rect 2658 5414 2710 5466
rect 2710 5414 2712 5466
rect 2736 5414 2774 5466
rect 2774 5414 2786 5466
rect 2786 5414 2792 5466
rect 2816 5414 2838 5466
rect 2838 5414 2850 5466
rect 2850 5414 2872 5466
rect 2896 5414 2902 5466
rect 2902 5414 2914 5466
rect 2914 5414 2952 5466
rect 2976 5414 2978 5466
rect 2978 5414 3030 5466
rect 3030 5414 3032 5466
rect 2656 5412 2712 5414
rect 2736 5412 2792 5414
rect 2816 5412 2872 5414
rect 2896 5412 2952 5414
rect 2976 5412 3032 5414
rect 1916 4922 1972 4924
rect 1996 4922 2052 4924
rect 2076 4922 2132 4924
rect 2156 4922 2212 4924
rect 2236 4922 2292 4924
rect 1916 4870 1918 4922
rect 1918 4870 1970 4922
rect 1970 4870 1972 4922
rect 1996 4870 2034 4922
rect 2034 4870 2046 4922
rect 2046 4870 2052 4922
rect 2076 4870 2098 4922
rect 2098 4870 2110 4922
rect 2110 4870 2132 4922
rect 2156 4870 2162 4922
rect 2162 4870 2174 4922
rect 2174 4870 2212 4922
rect 2236 4870 2238 4922
rect 2238 4870 2290 4922
rect 2290 4870 2292 4922
rect 1916 4868 1972 4870
rect 1996 4868 2052 4870
rect 2076 4868 2132 4870
rect 2156 4868 2212 4870
rect 2236 4868 2292 4870
rect 2656 4378 2712 4380
rect 2736 4378 2792 4380
rect 2816 4378 2872 4380
rect 2896 4378 2952 4380
rect 2976 4378 3032 4380
rect 2656 4326 2658 4378
rect 2658 4326 2710 4378
rect 2710 4326 2712 4378
rect 2736 4326 2774 4378
rect 2774 4326 2786 4378
rect 2786 4326 2792 4378
rect 2816 4326 2838 4378
rect 2838 4326 2850 4378
rect 2850 4326 2872 4378
rect 2896 4326 2902 4378
rect 2902 4326 2914 4378
rect 2914 4326 2952 4378
rect 2976 4326 2978 4378
rect 2978 4326 3030 4378
rect 3030 4326 3032 4378
rect 2656 4324 2712 4326
rect 2736 4324 2792 4326
rect 2816 4324 2872 4326
rect 2896 4324 2952 4326
rect 2976 4324 3032 4326
rect 3514 6160 3570 6216
rect 3606 5616 3662 5672
rect 5354 17720 5410 17776
rect 4802 15544 4858 15600
rect 5354 15952 5410 16008
rect 3790 7656 3846 7712
rect 3790 6432 3846 6488
rect 4342 7248 4398 7304
rect 4802 10648 4858 10704
rect 8656 23962 8712 23964
rect 8736 23962 8792 23964
rect 8816 23962 8872 23964
rect 8896 23962 8952 23964
rect 8976 23962 9032 23964
rect 8656 23910 8658 23962
rect 8658 23910 8710 23962
rect 8710 23910 8712 23962
rect 8736 23910 8774 23962
rect 8774 23910 8786 23962
rect 8786 23910 8792 23962
rect 8816 23910 8838 23962
rect 8838 23910 8850 23962
rect 8850 23910 8872 23962
rect 8896 23910 8902 23962
rect 8902 23910 8914 23962
rect 8914 23910 8952 23962
rect 8976 23910 8978 23962
rect 8978 23910 9030 23962
rect 9030 23910 9032 23962
rect 8656 23908 8712 23910
rect 8736 23908 8792 23910
rect 8816 23908 8872 23910
rect 8896 23908 8952 23910
rect 8976 23908 9032 23910
rect 7916 23418 7972 23420
rect 7996 23418 8052 23420
rect 8076 23418 8132 23420
rect 8156 23418 8212 23420
rect 8236 23418 8292 23420
rect 7916 23366 7918 23418
rect 7918 23366 7970 23418
rect 7970 23366 7972 23418
rect 7996 23366 8034 23418
rect 8034 23366 8046 23418
rect 8046 23366 8052 23418
rect 8076 23366 8098 23418
rect 8098 23366 8110 23418
rect 8110 23366 8132 23418
rect 8156 23366 8162 23418
rect 8162 23366 8174 23418
rect 8174 23366 8212 23418
rect 8236 23366 8238 23418
rect 8238 23366 8290 23418
rect 8290 23366 8292 23418
rect 7916 23364 7972 23366
rect 7996 23364 8052 23366
rect 8076 23364 8132 23366
rect 8156 23364 8212 23366
rect 8236 23364 8292 23366
rect 8656 22874 8712 22876
rect 8736 22874 8792 22876
rect 8816 22874 8872 22876
rect 8896 22874 8952 22876
rect 8976 22874 9032 22876
rect 8656 22822 8658 22874
rect 8658 22822 8710 22874
rect 8710 22822 8712 22874
rect 8736 22822 8774 22874
rect 8774 22822 8786 22874
rect 8786 22822 8792 22874
rect 8816 22822 8838 22874
rect 8838 22822 8850 22874
rect 8850 22822 8872 22874
rect 8896 22822 8902 22874
rect 8902 22822 8914 22874
rect 8914 22822 8952 22874
rect 8976 22822 8978 22874
rect 8978 22822 9030 22874
rect 9030 22822 9032 22874
rect 8656 22820 8712 22822
rect 8736 22820 8792 22822
rect 8816 22820 8872 22822
rect 8896 22820 8952 22822
rect 8976 22820 9032 22822
rect 7916 22330 7972 22332
rect 7996 22330 8052 22332
rect 8076 22330 8132 22332
rect 8156 22330 8212 22332
rect 8236 22330 8292 22332
rect 7916 22278 7918 22330
rect 7918 22278 7970 22330
rect 7970 22278 7972 22330
rect 7996 22278 8034 22330
rect 8034 22278 8046 22330
rect 8046 22278 8052 22330
rect 8076 22278 8098 22330
rect 8098 22278 8110 22330
rect 8110 22278 8132 22330
rect 8156 22278 8162 22330
rect 8162 22278 8174 22330
rect 8174 22278 8212 22330
rect 8236 22278 8238 22330
rect 8238 22278 8290 22330
rect 8290 22278 8292 22330
rect 7916 22276 7972 22278
rect 7996 22276 8052 22278
rect 8076 22276 8132 22278
rect 8156 22276 8212 22278
rect 8236 22276 8292 22278
rect 7916 21242 7972 21244
rect 7996 21242 8052 21244
rect 8076 21242 8132 21244
rect 8156 21242 8212 21244
rect 8236 21242 8292 21244
rect 7916 21190 7918 21242
rect 7918 21190 7970 21242
rect 7970 21190 7972 21242
rect 7996 21190 8034 21242
rect 8034 21190 8046 21242
rect 8046 21190 8052 21242
rect 8076 21190 8098 21242
rect 8098 21190 8110 21242
rect 8110 21190 8132 21242
rect 8156 21190 8162 21242
rect 8162 21190 8174 21242
rect 8174 21190 8212 21242
rect 8236 21190 8238 21242
rect 8238 21190 8290 21242
rect 8290 21190 8292 21242
rect 7916 21188 7972 21190
rect 7996 21188 8052 21190
rect 8076 21188 8132 21190
rect 8156 21188 8212 21190
rect 8236 21188 8292 21190
rect 7916 20154 7972 20156
rect 7996 20154 8052 20156
rect 8076 20154 8132 20156
rect 8156 20154 8212 20156
rect 8236 20154 8292 20156
rect 7916 20102 7918 20154
rect 7918 20102 7970 20154
rect 7970 20102 7972 20154
rect 7996 20102 8034 20154
rect 8034 20102 8046 20154
rect 8046 20102 8052 20154
rect 8076 20102 8098 20154
rect 8098 20102 8110 20154
rect 8110 20102 8132 20154
rect 8156 20102 8162 20154
rect 8162 20102 8174 20154
rect 8174 20102 8212 20154
rect 8236 20102 8238 20154
rect 8238 20102 8290 20154
rect 8290 20102 8292 20154
rect 7916 20100 7972 20102
rect 7996 20100 8052 20102
rect 8076 20100 8132 20102
rect 8156 20100 8212 20102
rect 8236 20100 8292 20102
rect 8656 21786 8712 21788
rect 8736 21786 8792 21788
rect 8816 21786 8872 21788
rect 8896 21786 8952 21788
rect 8976 21786 9032 21788
rect 8656 21734 8658 21786
rect 8658 21734 8710 21786
rect 8710 21734 8712 21786
rect 8736 21734 8774 21786
rect 8774 21734 8786 21786
rect 8786 21734 8792 21786
rect 8816 21734 8838 21786
rect 8838 21734 8850 21786
rect 8850 21734 8872 21786
rect 8896 21734 8902 21786
rect 8902 21734 8914 21786
rect 8914 21734 8952 21786
rect 8976 21734 8978 21786
rect 8978 21734 9030 21786
rect 9030 21734 9032 21786
rect 8656 21732 8712 21734
rect 8736 21732 8792 21734
rect 8816 21732 8872 21734
rect 8896 21732 8952 21734
rect 8976 21732 9032 21734
rect 8656 20698 8712 20700
rect 8736 20698 8792 20700
rect 8816 20698 8872 20700
rect 8896 20698 8952 20700
rect 8976 20698 9032 20700
rect 8656 20646 8658 20698
rect 8658 20646 8710 20698
rect 8710 20646 8712 20698
rect 8736 20646 8774 20698
rect 8774 20646 8786 20698
rect 8786 20646 8792 20698
rect 8816 20646 8838 20698
rect 8838 20646 8850 20698
rect 8850 20646 8872 20698
rect 8896 20646 8902 20698
rect 8902 20646 8914 20698
rect 8914 20646 8952 20698
rect 8976 20646 8978 20698
rect 8978 20646 9030 20698
rect 9030 20646 9032 20698
rect 8656 20644 8712 20646
rect 8736 20644 8792 20646
rect 8816 20644 8872 20646
rect 8896 20644 8952 20646
rect 8976 20644 9032 20646
rect 7916 19066 7972 19068
rect 7996 19066 8052 19068
rect 8076 19066 8132 19068
rect 8156 19066 8212 19068
rect 8236 19066 8292 19068
rect 7916 19014 7918 19066
rect 7918 19014 7970 19066
rect 7970 19014 7972 19066
rect 7996 19014 8034 19066
rect 8034 19014 8046 19066
rect 8046 19014 8052 19066
rect 8076 19014 8098 19066
rect 8098 19014 8110 19066
rect 8110 19014 8132 19066
rect 8156 19014 8162 19066
rect 8162 19014 8174 19066
rect 8174 19014 8212 19066
rect 8236 19014 8238 19066
rect 8238 19014 8290 19066
rect 8290 19014 8292 19066
rect 7916 19012 7972 19014
rect 7996 19012 8052 19014
rect 8076 19012 8132 19014
rect 8156 19012 8212 19014
rect 8236 19012 8292 19014
rect 3974 6568 4030 6624
rect 3974 5888 4030 5944
rect 4526 6840 4582 6896
rect 4618 6704 4674 6760
rect 4802 7656 4858 7712
rect 1916 3834 1972 3836
rect 1996 3834 2052 3836
rect 2076 3834 2132 3836
rect 2156 3834 2212 3836
rect 2236 3834 2292 3836
rect 1916 3782 1918 3834
rect 1918 3782 1970 3834
rect 1970 3782 1972 3834
rect 1996 3782 2034 3834
rect 2034 3782 2046 3834
rect 2046 3782 2052 3834
rect 2076 3782 2098 3834
rect 2098 3782 2110 3834
rect 2110 3782 2132 3834
rect 2156 3782 2162 3834
rect 2162 3782 2174 3834
rect 2174 3782 2212 3834
rect 2236 3782 2238 3834
rect 2238 3782 2290 3834
rect 2290 3782 2292 3834
rect 1916 3780 1972 3782
rect 1996 3780 2052 3782
rect 2076 3780 2132 3782
rect 2156 3780 2212 3782
rect 2236 3780 2292 3782
rect 2656 3290 2712 3292
rect 2736 3290 2792 3292
rect 2816 3290 2872 3292
rect 2896 3290 2952 3292
rect 2976 3290 3032 3292
rect 2656 3238 2658 3290
rect 2658 3238 2710 3290
rect 2710 3238 2712 3290
rect 2736 3238 2774 3290
rect 2774 3238 2786 3290
rect 2786 3238 2792 3290
rect 2816 3238 2838 3290
rect 2838 3238 2850 3290
rect 2850 3238 2872 3290
rect 2896 3238 2902 3290
rect 2902 3238 2914 3290
rect 2914 3238 2952 3290
rect 2976 3238 2978 3290
rect 2978 3238 3030 3290
rect 3030 3238 3032 3290
rect 2656 3236 2712 3238
rect 2736 3236 2792 3238
rect 2816 3236 2872 3238
rect 2896 3236 2952 3238
rect 2976 3236 3032 3238
rect 5446 7112 5502 7168
rect 5354 6976 5410 7032
rect 1916 2746 1972 2748
rect 1996 2746 2052 2748
rect 2076 2746 2132 2748
rect 2156 2746 2212 2748
rect 2236 2746 2292 2748
rect 1916 2694 1918 2746
rect 1918 2694 1970 2746
rect 1970 2694 1972 2746
rect 1996 2694 2034 2746
rect 2034 2694 2046 2746
rect 2046 2694 2052 2746
rect 2076 2694 2098 2746
rect 2098 2694 2110 2746
rect 2110 2694 2132 2746
rect 2156 2694 2162 2746
rect 2162 2694 2174 2746
rect 2174 2694 2212 2746
rect 2236 2694 2238 2746
rect 2238 2694 2290 2746
rect 2290 2694 2292 2746
rect 1916 2692 1972 2694
rect 1996 2692 2052 2694
rect 2076 2692 2132 2694
rect 2156 2692 2212 2694
rect 2236 2692 2292 2694
rect 6458 9560 6514 9616
rect 7102 7928 7158 7984
rect 7916 17978 7972 17980
rect 7996 17978 8052 17980
rect 8076 17978 8132 17980
rect 8156 17978 8212 17980
rect 8236 17978 8292 17980
rect 7916 17926 7918 17978
rect 7918 17926 7970 17978
rect 7970 17926 7972 17978
rect 7996 17926 8034 17978
rect 8034 17926 8046 17978
rect 8046 17926 8052 17978
rect 8076 17926 8098 17978
rect 8098 17926 8110 17978
rect 8110 17926 8132 17978
rect 8156 17926 8162 17978
rect 8162 17926 8174 17978
rect 8174 17926 8212 17978
rect 8236 17926 8238 17978
rect 8238 17926 8290 17978
rect 8290 17926 8292 17978
rect 7916 17924 7972 17926
rect 7996 17924 8052 17926
rect 8076 17924 8132 17926
rect 8156 17924 8212 17926
rect 8236 17924 8292 17926
rect 7916 16890 7972 16892
rect 7996 16890 8052 16892
rect 8076 16890 8132 16892
rect 8156 16890 8212 16892
rect 8236 16890 8292 16892
rect 7916 16838 7918 16890
rect 7918 16838 7970 16890
rect 7970 16838 7972 16890
rect 7996 16838 8034 16890
rect 8034 16838 8046 16890
rect 8046 16838 8052 16890
rect 8076 16838 8098 16890
rect 8098 16838 8110 16890
rect 8110 16838 8132 16890
rect 8156 16838 8162 16890
rect 8162 16838 8174 16890
rect 8174 16838 8212 16890
rect 8236 16838 8238 16890
rect 8238 16838 8290 16890
rect 8290 16838 8292 16890
rect 7916 16836 7972 16838
rect 7996 16836 8052 16838
rect 8076 16836 8132 16838
rect 8156 16836 8212 16838
rect 8236 16836 8292 16838
rect 8298 15952 8354 16008
rect 7916 15802 7972 15804
rect 7996 15802 8052 15804
rect 8076 15802 8132 15804
rect 8156 15802 8212 15804
rect 8236 15802 8292 15804
rect 7916 15750 7918 15802
rect 7918 15750 7970 15802
rect 7970 15750 7972 15802
rect 7996 15750 8034 15802
rect 8034 15750 8046 15802
rect 8046 15750 8052 15802
rect 8076 15750 8098 15802
rect 8098 15750 8110 15802
rect 8110 15750 8132 15802
rect 8156 15750 8162 15802
rect 8162 15750 8174 15802
rect 8174 15750 8212 15802
rect 8236 15750 8238 15802
rect 8238 15750 8290 15802
rect 8290 15750 8292 15802
rect 7916 15748 7972 15750
rect 7996 15748 8052 15750
rect 8076 15748 8132 15750
rect 8156 15748 8212 15750
rect 8236 15748 8292 15750
rect 8656 19610 8712 19612
rect 8736 19610 8792 19612
rect 8816 19610 8872 19612
rect 8896 19610 8952 19612
rect 8976 19610 9032 19612
rect 8656 19558 8658 19610
rect 8658 19558 8710 19610
rect 8710 19558 8712 19610
rect 8736 19558 8774 19610
rect 8774 19558 8786 19610
rect 8786 19558 8792 19610
rect 8816 19558 8838 19610
rect 8838 19558 8850 19610
rect 8850 19558 8872 19610
rect 8896 19558 8902 19610
rect 8902 19558 8914 19610
rect 8914 19558 8952 19610
rect 8976 19558 8978 19610
rect 8978 19558 9030 19610
rect 9030 19558 9032 19610
rect 8656 19556 8712 19558
rect 8736 19556 8792 19558
rect 8816 19556 8872 19558
rect 8896 19556 8952 19558
rect 8976 19556 9032 19558
rect 8656 18522 8712 18524
rect 8736 18522 8792 18524
rect 8816 18522 8872 18524
rect 8896 18522 8952 18524
rect 8976 18522 9032 18524
rect 8656 18470 8658 18522
rect 8658 18470 8710 18522
rect 8710 18470 8712 18522
rect 8736 18470 8774 18522
rect 8774 18470 8786 18522
rect 8786 18470 8792 18522
rect 8816 18470 8838 18522
rect 8838 18470 8850 18522
rect 8850 18470 8872 18522
rect 8896 18470 8902 18522
rect 8902 18470 8914 18522
rect 8914 18470 8952 18522
rect 8976 18470 8978 18522
rect 8978 18470 9030 18522
rect 9030 18470 9032 18522
rect 8656 18468 8712 18470
rect 8736 18468 8792 18470
rect 8816 18468 8872 18470
rect 8896 18468 8952 18470
rect 8976 18468 9032 18470
rect 8656 17434 8712 17436
rect 8736 17434 8792 17436
rect 8816 17434 8872 17436
rect 8896 17434 8952 17436
rect 8976 17434 9032 17436
rect 8656 17382 8658 17434
rect 8658 17382 8710 17434
rect 8710 17382 8712 17434
rect 8736 17382 8774 17434
rect 8774 17382 8786 17434
rect 8786 17382 8792 17434
rect 8816 17382 8838 17434
rect 8838 17382 8850 17434
rect 8850 17382 8872 17434
rect 8896 17382 8902 17434
rect 8902 17382 8914 17434
rect 8914 17382 8952 17434
rect 8976 17382 8978 17434
rect 8978 17382 9030 17434
rect 9030 17382 9032 17434
rect 8656 17380 8712 17382
rect 8736 17380 8792 17382
rect 8816 17380 8872 17382
rect 8896 17380 8952 17382
rect 8976 17380 9032 17382
rect 8666 17040 8722 17096
rect 9034 16668 9036 16688
rect 9036 16668 9088 16688
rect 9088 16668 9090 16688
rect 9034 16632 9090 16668
rect 8656 16346 8712 16348
rect 8736 16346 8792 16348
rect 8816 16346 8872 16348
rect 8896 16346 8952 16348
rect 8976 16346 9032 16348
rect 8656 16294 8658 16346
rect 8658 16294 8710 16346
rect 8710 16294 8712 16346
rect 8736 16294 8774 16346
rect 8774 16294 8786 16346
rect 8786 16294 8792 16346
rect 8816 16294 8838 16346
rect 8838 16294 8850 16346
rect 8850 16294 8872 16346
rect 8896 16294 8902 16346
rect 8902 16294 8914 16346
rect 8914 16294 8952 16346
rect 8976 16294 8978 16346
rect 8978 16294 9030 16346
rect 9030 16294 9032 16346
rect 8656 16292 8712 16294
rect 8736 16292 8792 16294
rect 8816 16292 8872 16294
rect 8896 16292 8952 16294
rect 8976 16292 9032 16294
rect 9126 16088 9182 16144
rect 8656 15258 8712 15260
rect 8736 15258 8792 15260
rect 8816 15258 8872 15260
rect 8896 15258 8952 15260
rect 8976 15258 9032 15260
rect 8656 15206 8658 15258
rect 8658 15206 8710 15258
rect 8710 15206 8712 15258
rect 8736 15206 8774 15258
rect 8774 15206 8786 15258
rect 8786 15206 8792 15258
rect 8816 15206 8838 15258
rect 8838 15206 8850 15258
rect 8850 15206 8872 15258
rect 8896 15206 8902 15258
rect 8902 15206 8914 15258
rect 8914 15206 8952 15258
rect 8976 15206 8978 15258
rect 8978 15206 9030 15258
rect 9030 15206 9032 15258
rect 8656 15204 8712 15206
rect 8736 15204 8792 15206
rect 8816 15204 8872 15206
rect 8896 15204 8952 15206
rect 8976 15204 9032 15206
rect 7916 14714 7972 14716
rect 7996 14714 8052 14716
rect 8076 14714 8132 14716
rect 8156 14714 8212 14716
rect 8236 14714 8292 14716
rect 7916 14662 7918 14714
rect 7918 14662 7970 14714
rect 7970 14662 7972 14714
rect 7996 14662 8034 14714
rect 8034 14662 8046 14714
rect 8046 14662 8052 14714
rect 8076 14662 8098 14714
rect 8098 14662 8110 14714
rect 8110 14662 8132 14714
rect 8156 14662 8162 14714
rect 8162 14662 8174 14714
rect 8174 14662 8212 14714
rect 8236 14662 8238 14714
rect 8238 14662 8290 14714
rect 8290 14662 8292 14714
rect 7916 14660 7972 14662
rect 7996 14660 8052 14662
rect 8076 14660 8132 14662
rect 8156 14660 8212 14662
rect 8236 14660 8292 14662
rect 7916 13626 7972 13628
rect 7996 13626 8052 13628
rect 8076 13626 8132 13628
rect 8156 13626 8212 13628
rect 8236 13626 8292 13628
rect 7916 13574 7918 13626
rect 7918 13574 7970 13626
rect 7970 13574 7972 13626
rect 7996 13574 8034 13626
rect 8034 13574 8046 13626
rect 8046 13574 8052 13626
rect 8076 13574 8098 13626
rect 8098 13574 8110 13626
rect 8110 13574 8132 13626
rect 8156 13574 8162 13626
rect 8162 13574 8174 13626
rect 8174 13574 8212 13626
rect 8236 13574 8238 13626
rect 8238 13574 8290 13626
rect 8290 13574 8292 13626
rect 7916 13572 7972 13574
rect 7996 13572 8052 13574
rect 8076 13572 8132 13574
rect 8156 13572 8212 13574
rect 8236 13572 8292 13574
rect 8656 14170 8712 14172
rect 8736 14170 8792 14172
rect 8816 14170 8872 14172
rect 8896 14170 8952 14172
rect 8976 14170 9032 14172
rect 8656 14118 8658 14170
rect 8658 14118 8710 14170
rect 8710 14118 8712 14170
rect 8736 14118 8774 14170
rect 8774 14118 8786 14170
rect 8786 14118 8792 14170
rect 8816 14118 8838 14170
rect 8838 14118 8850 14170
rect 8850 14118 8872 14170
rect 8896 14118 8902 14170
rect 8902 14118 8914 14170
rect 8914 14118 8952 14170
rect 8976 14118 8978 14170
rect 8978 14118 9030 14170
rect 9030 14118 9032 14170
rect 8656 14116 8712 14118
rect 8736 14116 8792 14118
rect 8816 14116 8872 14118
rect 8896 14116 8952 14118
rect 8976 14116 9032 14118
rect 8656 13082 8712 13084
rect 8736 13082 8792 13084
rect 8816 13082 8872 13084
rect 8896 13082 8952 13084
rect 8976 13082 9032 13084
rect 8656 13030 8658 13082
rect 8658 13030 8710 13082
rect 8710 13030 8712 13082
rect 8736 13030 8774 13082
rect 8774 13030 8786 13082
rect 8786 13030 8792 13082
rect 8816 13030 8838 13082
rect 8838 13030 8850 13082
rect 8850 13030 8872 13082
rect 8896 13030 8902 13082
rect 8902 13030 8914 13082
rect 8914 13030 8952 13082
rect 8976 13030 8978 13082
rect 8978 13030 9030 13082
rect 9030 13030 9032 13082
rect 8656 13028 8712 13030
rect 8736 13028 8792 13030
rect 8816 13028 8872 13030
rect 8896 13028 8952 13030
rect 8976 13028 9032 13030
rect 8390 12844 8446 12880
rect 8390 12824 8392 12844
rect 8392 12824 8444 12844
rect 8444 12824 8446 12844
rect 7916 12538 7972 12540
rect 7996 12538 8052 12540
rect 8076 12538 8132 12540
rect 8156 12538 8212 12540
rect 8236 12538 8292 12540
rect 7916 12486 7918 12538
rect 7918 12486 7970 12538
rect 7970 12486 7972 12538
rect 7996 12486 8034 12538
rect 8034 12486 8046 12538
rect 8046 12486 8052 12538
rect 8076 12486 8098 12538
rect 8098 12486 8110 12538
rect 8110 12486 8132 12538
rect 8156 12486 8162 12538
rect 8162 12486 8174 12538
rect 8174 12486 8212 12538
rect 8236 12486 8238 12538
rect 8238 12486 8290 12538
rect 8290 12486 8292 12538
rect 7916 12484 7972 12486
rect 7996 12484 8052 12486
rect 8076 12484 8132 12486
rect 8156 12484 8212 12486
rect 8236 12484 8292 12486
rect 7916 11450 7972 11452
rect 7996 11450 8052 11452
rect 8076 11450 8132 11452
rect 8156 11450 8212 11452
rect 8236 11450 8292 11452
rect 7916 11398 7918 11450
rect 7918 11398 7970 11450
rect 7970 11398 7972 11450
rect 7996 11398 8034 11450
rect 8034 11398 8046 11450
rect 8046 11398 8052 11450
rect 8076 11398 8098 11450
rect 8098 11398 8110 11450
rect 8110 11398 8132 11450
rect 8156 11398 8162 11450
rect 8162 11398 8174 11450
rect 8174 11398 8212 11450
rect 8236 11398 8238 11450
rect 8238 11398 8290 11450
rect 8290 11398 8292 11450
rect 7916 11396 7972 11398
rect 7996 11396 8052 11398
rect 8076 11396 8132 11398
rect 8156 11396 8212 11398
rect 8236 11396 8292 11398
rect 7916 10362 7972 10364
rect 7996 10362 8052 10364
rect 8076 10362 8132 10364
rect 8156 10362 8212 10364
rect 8236 10362 8292 10364
rect 7916 10310 7918 10362
rect 7918 10310 7970 10362
rect 7970 10310 7972 10362
rect 7996 10310 8034 10362
rect 8034 10310 8046 10362
rect 8046 10310 8052 10362
rect 8076 10310 8098 10362
rect 8098 10310 8110 10362
rect 8110 10310 8132 10362
rect 8156 10310 8162 10362
rect 8162 10310 8174 10362
rect 8174 10310 8212 10362
rect 8236 10310 8238 10362
rect 8238 10310 8290 10362
rect 8290 10310 8292 10362
rect 7916 10308 7972 10310
rect 7996 10308 8052 10310
rect 8076 10308 8132 10310
rect 8156 10308 8212 10310
rect 8236 10308 8292 10310
rect 7916 9274 7972 9276
rect 7996 9274 8052 9276
rect 8076 9274 8132 9276
rect 8156 9274 8212 9276
rect 8236 9274 8292 9276
rect 7916 9222 7918 9274
rect 7918 9222 7970 9274
rect 7970 9222 7972 9274
rect 7996 9222 8034 9274
rect 8034 9222 8046 9274
rect 8046 9222 8052 9274
rect 8076 9222 8098 9274
rect 8098 9222 8110 9274
rect 8110 9222 8132 9274
rect 8156 9222 8162 9274
rect 8162 9222 8174 9274
rect 8174 9222 8212 9274
rect 8236 9222 8238 9274
rect 8238 9222 8290 9274
rect 8290 9222 8292 9274
rect 7916 9220 7972 9222
rect 7996 9220 8052 9222
rect 8076 9220 8132 9222
rect 8156 9220 8212 9222
rect 8236 9220 8292 9222
rect 8656 11994 8712 11996
rect 8736 11994 8792 11996
rect 8816 11994 8872 11996
rect 8896 11994 8952 11996
rect 8976 11994 9032 11996
rect 8656 11942 8658 11994
rect 8658 11942 8710 11994
rect 8710 11942 8712 11994
rect 8736 11942 8774 11994
rect 8774 11942 8786 11994
rect 8786 11942 8792 11994
rect 8816 11942 8838 11994
rect 8838 11942 8850 11994
rect 8850 11942 8872 11994
rect 8896 11942 8902 11994
rect 8902 11942 8914 11994
rect 8914 11942 8952 11994
rect 8976 11942 8978 11994
rect 8978 11942 9030 11994
rect 9030 11942 9032 11994
rect 8656 11940 8712 11942
rect 8736 11940 8792 11942
rect 8816 11940 8872 11942
rect 8896 11940 8952 11942
rect 8976 11940 9032 11942
rect 10138 17720 10194 17776
rect 9402 12688 9458 12744
rect 9402 12588 9404 12608
rect 9404 12588 9456 12608
rect 9456 12588 9458 12608
rect 9402 12552 9458 12588
rect 8656 10906 8712 10908
rect 8736 10906 8792 10908
rect 8816 10906 8872 10908
rect 8896 10906 8952 10908
rect 8976 10906 9032 10908
rect 8656 10854 8658 10906
rect 8658 10854 8710 10906
rect 8710 10854 8712 10906
rect 8736 10854 8774 10906
rect 8774 10854 8786 10906
rect 8786 10854 8792 10906
rect 8816 10854 8838 10906
rect 8838 10854 8850 10906
rect 8850 10854 8872 10906
rect 8896 10854 8902 10906
rect 8902 10854 8914 10906
rect 8914 10854 8952 10906
rect 8976 10854 8978 10906
rect 8978 10854 9030 10906
rect 9030 10854 9032 10906
rect 8656 10852 8712 10854
rect 8736 10852 8792 10854
rect 8816 10852 8872 10854
rect 8896 10852 8952 10854
rect 8976 10852 9032 10854
rect 8656 9818 8712 9820
rect 8736 9818 8792 9820
rect 8816 9818 8872 9820
rect 8896 9818 8952 9820
rect 8976 9818 9032 9820
rect 8656 9766 8658 9818
rect 8658 9766 8710 9818
rect 8710 9766 8712 9818
rect 8736 9766 8774 9818
rect 8774 9766 8786 9818
rect 8786 9766 8792 9818
rect 8816 9766 8838 9818
rect 8838 9766 8850 9818
rect 8850 9766 8872 9818
rect 8896 9766 8902 9818
rect 8902 9766 8914 9818
rect 8914 9766 8952 9818
rect 8976 9766 8978 9818
rect 8978 9766 9030 9818
rect 9030 9766 9032 9818
rect 8656 9764 8712 9766
rect 8736 9764 8792 9766
rect 8816 9764 8872 9766
rect 8896 9764 8952 9766
rect 8976 9764 9032 9766
rect 7916 8186 7972 8188
rect 7996 8186 8052 8188
rect 8076 8186 8132 8188
rect 8156 8186 8212 8188
rect 8236 8186 8292 8188
rect 7916 8134 7918 8186
rect 7918 8134 7970 8186
rect 7970 8134 7972 8186
rect 7996 8134 8034 8186
rect 8034 8134 8046 8186
rect 8046 8134 8052 8186
rect 8076 8134 8098 8186
rect 8098 8134 8110 8186
rect 8110 8134 8132 8186
rect 8156 8134 8162 8186
rect 8162 8134 8174 8186
rect 8174 8134 8212 8186
rect 8236 8134 8238 8186
rect 8238 8134 8290 8186
rect 8290 8134 8292 8186
rect 7916 8132 7972 8134
rect 7996 8132 8052 8134
rect 8076 8132 8132 8134
rect 8156 8132 8212 8134
rect 8236 8132 8292 8134
rect 8656 8730 8712 8732
rect 8736 8730 8792 8732
rect 8816 8730 8872 8732
rect 8896 8730 8952 8732
rect 8976 8730 9032 8732
rect 8656 8678 8658 8730
rect 8658 8678 8710 8730
rect 8710 8678 8712 8730
rect 8736 8678 8774 8730
rect 8774 8678 8786 8730
rect 8786 8678 8792 8730
rect 8816 8678 8838 8730
rect 8838 8678 8850 8730
rect 8850 8678 8872 8730
rect 8896 8678 8902 8730
rect 8902 8678 8914 8730
rect 8914 8678 8952 8730
rect 8976 8678 8978 8730
rect 8978 8678 9030 8730
rect 9030 8678 9032 8730
rect 8656 8676 8712 8678
rect 8736 8676 8792 8678
rect 8816 8676 8872 8678
rect 8896 8676 8952 8678
rect 8976 8676 9032 8678
rect 7010 6704 7066 6760
rect 6918 6452 6974 6488
rect 6918 6432 6920 6452
rect 6920 6432 6972 6452
rect 6972 6432 6974 6452
rect 6734 6296 6790 6352
rect 6458 5752 6514 5808
rect 8574 7792 8630 7848
rect 7916 7098 7972 7100
rect 7996 7098 8052 7100
rect 8076 7098 8132 7100
rect 8156 7098 8212 7100
rect 8236 7098 8292 7100
rect 7916 7046 7918 7098
rect 7918 7046 7970 7098
rect 7970 7046 7972 7098
rect 7996 7046 8034 7098
rect 8034 7046 8046 7098
rect 8046 7046 8052 7098
rect 8076 7046 8098 7098
rect 8098 7046 8110 7098
rect 8110 7046 8132 7098
rect 8156 7046 8162 7098
rect 8162 7046 8174 7098
rect 8174 7046 8212 7098
rect 8236 7046 8238 7098
rect 8238 7046 8290 7098
rect 8290 7046 8292 7098
rect 7916 7044 7972 7046
rect 7996 7044 8052 7046
rect 8076 7044 8132 7046
rect 8156 7044 8212 7046
rect 8236 7044 8292 7046
rect 8298 6160 8354 6216
rect 7916 6010 7972 6012
rect 7996 6010 8052 6012
rect 8076 6010 8132 6012
rect 8156 6010 8212 6012
rect 8236 6010 8292 6012
rect 7916 5958 7918 6010
rect 7918 5958 7970 6010
rect 7970 5958 7972 6010
rect 7996 5958 8034 6010
rect 8034 5958 8046 6010
rect 8046 5958 8052 6010
rect 8076 5958 8098 6010
rect 8098 5958 8110 6010
rect 8110 5958 8132 6010
rect 8156 5958 8162 6010
rect 8162 5958 8174 6010
rect 8174 5958 8212 6010
rect 8236 5958 8238 6010
rect 8238 5958 8290 6010
rect 8290 5958 8292 6010
rect 7916 5956 7972 5958
rect 7996 5956 8052 5958
rect 8076 5956 8132 5958
rect 8156 5956 8212 5958
rect 8236 5956 8292 5958
rect 7916 4922 7972 4924
rect 7996 4922 8052 4924
rect 8076 4922 8132 4924
rect 8156 4922 8212 4924
rect 8236 4922 8292 4924
rect 7916 4870 7918 4922
rect 7918 4870 7970 4922
rect 7970 4870 7972 4922
rect 7996 4870 8034 4922
rect 8034 4870 8046 4922
rect 8046 4870 8052 4922
rect 8076 4870 8098 4922
rect 8098 4870 8110 4922
rect 8110 4870 8132 4922
rect 8156 4870 8162 4922
rect 8162 4870 8174 4922
rect 8174 4870 8212 4922
rect 8236 4870 8238 4922
rect 8238 4870 8290 4922
rect 8290 4870 8292 4922
rect 7916 4868 7972 4870
rect 7996 4868 8052 4870
rect 8076 4868 8132 4870
rect 8156 4868 8212 4870
rect 8236 4868 8292 4870
rect 7916 3834 7972 3836
rect 7996 3834 8052 3836
rect 8076 3834 8132 3836
rect 8156 3834 8212 3836
rect 8236 3834 8292 3836
rect 7916 3782 7918 3834
rect 7918 3782 7970 3834
rect 7970 3782 7972 3834
rect 7996 3782 8034 3834
rect 8034 3782 8046 3834
rect 8046 3782 8052 3834
rect 8076 3782 8098 3834
rect 8098 3782 8110 3834
rect 8110 3782 8132 3834
rect 8156 3782 8162 3834
rect 8162 3782 8174 3834
rect 8174 3782 8212 3834
rect 8236 3782 8238 3834
rect 8238 3782 8290 3834
rect 8290 3782 8292 3834
rect 7916 3780 7972 3782
rect 7996 3780 8052 3782
rect 8076 3780 8132 3782
rect 8156 3780 8212 3782
rect 8236 3780 8292 3782
rect 8656 7642 8712 7644
rect 8736 7642 8792 7644
rect 8816 7642 8872 7644
rect 8896 7642 8952 7644
rect 8976 7642 9032 7644
rect 8656 7590 8658 7642
rect 8658 7590 8710 7642
rect 8710 7590 8712 7642
rect 8736 7590 8774 7642
rect 8774 7590 8786 7642
rect 8786 7590 8792 7642
rect 8816 7590 8838 7642
rect 8838 7590 8850 7642
rect 8850 7590 8872 7642
rect 8896 7590 8902 7642
rect 8902 7590 8914 7642
rect 8914 7590 8952 7642
rect 8976 7590 8978 7642
rect 8978 7590 9030 7642
rect 9030 7590 9032 7642
rect 8656 7588 8712 7590
rect 8736 7588 8792 7590
rect 8816 7588 8872 7590
rect 8896 7588 8952 7590
rect 8976 7588 9032 7590
rect 8656 6554 8712 6556
rect 8736 6554 8792 6556
rect 8816 6554 8872 6556
rect 8896 6554 8952 6556
rect 8976 6554 9032 6556
rect 8656 6502 8658 6554
rect 8658 6502 8710 6554
rect 8710 6502 8712 6554
rect 8736 6502 8774 6554
rect 8774 6502 8786 6554
rect 8786 6502 8792 6554
rect 8816 6502 8838 6554
rect 8838 6502 8850 6554
rect 8850 6502 8872 6554
rect 8896 6502 8902 6554
rect 8902 6502 8914 6554
rect 8914 6502 8952 6554
rect 8976 6502 8978 6554
rect 8978 6502 9030 6554
rect 9030 6502 9032 6554
rect 8656 6500 8712 6502
rect 8736 6500 8792 6502
rect 8816 6500 8872 6502
rect 8896 6500 8952 6502
rect 8976 6500 9032 6502
rect 9310 10648 9366 10704
rect 8656 5466 8712 5468
rect 8736 5466 8792 5468
rect 8816 5466 8872 5468
rect 8896 5466 8952 5468
rect 8976 5466 9032 5468
rect 8656 5414 8658 5466
rect 8658 5414 8710 5466
rect 8710 5414 8712 5466
rect 8736 5414 8774 5466
rect 8774 5414 8786 5466
rect 8786 5414 8792 5466
rect 8816 5414 8838 5466
rect 8838 5414 8850 5466
rect 8850 5414 8872 5466
rect 8896 5414 8902 5466
rect 8902 5414 8914 5466
rect 8914 5414 8952 5466
rect 8976 5414 8978 5466
rect 8978 5414 9030 5466
rect 9030 5414 9032 5466
rect 8656 5412 8712 5414
rect 8736 5412 8792 5414
rect 8816 5412 8872 5414
rect 8896 5412 8952 5414
rect 8976 5412 9032 5414
rect 8656 4378 8712 4380
rect 8736 4378 8792 4380
rect 8816 4378 8872 4380
rect 8896 4378 8952 4380
rect 8976 4378 9032 4380
rect 8656 4326 8658 4378
rect 8658 4326 8710 4378
rect 8710 4326 8712 4378
rect 8736 4326 8774 4378
rect 8774 4326 8786 4378
rect 8786 4326 8792 4378
rect 8816 4326 8838 4378
rect 8838 4326 8850 4378
rect 8850 4326 8872 4378
rect 8896 4326 8902 4378
rect 8902 4326 8914 4378
rect 8914 4326 8952 4378
rect 8976 4326 8978 4378
rect 8978 4326 9030 4378
rect 9030 4326 9032 4378
rect 8656 4324 8712 4326
rect 8736 4324 8792 4326
rect 8816 4324 8872 4326
rect 8896 4324 8952 4326
rect 8976 4324 9032 4326
rect 9770 12552 9826 12608
rect 13916 23418 13972 23420
rect 13996 23418 14052 23420
rect 14076 23418 14132 23420
rect 14156 23418 14212 23420
rect 14236 23418 14292 23420
rect 13916 23366 13918 23418
rect 13918 23366 13970 23418
rect 13970 23366 13972 23418
rect 13996 23366 14034 23418
rect 14034 23366 14046 23418
rect 14046 23366 14052 23418
rect 14076 23366 14098 23418
rect 14098 23366 14110 23418
rect 14110 23366 14132 23418
rect 14156 23366 14162 23418
rect 14162 23366 14174 23418
rect 14174 23366 14212 23418
rect 14236 23366 14238 23418
rect 14238 23366 14290 23418
rect 14290 23366 14292 23418
rect 13916 23364 13972 23366
rect 13996 23364 14052 23366
rect 14076 23364 14132 23366
rect 14156 23364 14212 23366
rect 14236 23364 14292 23366
rect 13916 22330 13972 22332
rect 13996 22330 14052 22332
rect 14076 22330 14132 22332
rect 14156 22330 14212 22332
rect 14236 22330 14292 22332
rect 13916 22278 13918 22330
rect 13918 22278 13970 22330
rect 13970 22278 13972 22330
rect 13996 22278 14034 22330
rect 14034 22278 14046 22330
rect 14046 22278 14052 22330
rect 14076 22278 14098 22330
rect 14098 22278 14110 22330
rect 14110 22278 14132 22330
rect 14156 22278 14162 22330
rect 14162 22278 14174 22330
rect 14174 22278 14212 22330
rect 14236 22278 14238 22330
rect 14238 22278 14290 22330
rect 14290 22278 14292 22330
rect 13916 22276 13972 22278
rect 13996 22276 14052 22278
rect 14076 22276 14132 22278
rect 14156 22276 14212 22278
rect 14236 22276 14292 22278
rect 13916 21242 13972 21244
rect 13996 21242 14052 21244
rect 14076 21242 14132 21244
rect 14156 21242 14212 21244
rect 14236 21242 14292 21244
rect 13916 21190 13918 21242
rect 13918 21190 13970 21242
rect 13970 21190 13972 21242
rect 13996 21190 14034 21242
rect 14034 21190 14046 21242
rect 14046 21190 14052 21242
rect 14076 21190 14098 21242
rect 14098 21190 14110 21242
rect 14110 21190 14132 21242
rect 14156 21190 14162 21242
rect 14162 21190 14174 21242
rect 14174 21190 14212 21242
rect 14236 21190 14238 21242
rect 14238 21190 14290 21242
rect 14290 21190 14292 21242
rect 13916 21188 13972 21190
rect 13996 21188 14052 21190
rect 14076 21188 14132 21190
rect 14156 21188 14212 21190
rect 14236 21188 14292 21190
rect 13916 20154 13972 20156
rect 13996 20154 14052 20156
rect 14076 20154 14132 20156
rect 14156 20154 14212 20156
rect 14236 20154 14292 20156
rect 13916 20102 13918 20154
rect 13918 20102 13970 20154
rect 13970 20102 13972 20154
rect 13996 20102 14034 20154
rect 14034 20102 14046 20154
rect 14046 20102 14052 20154
rect 14076 20102 14098 20154
rect 14098 20102 14110 20154
rect 14110 20102 14132 20154
rect 14156 20102 14162 20154
rect 14162 20102 14174 20154
rect 14174 20102 14212 20154
rect 14236 20102 14238 20154
rect 14238 20102 14290 20154
rect 14290 20102 14292 20154
rect 13916 20100 13972 20102
rect 13996 20100 14052 20102
rect 14076 20100 14132 20102
rect 14156 20100 14212 20102
rect 14236 20100 14292 20102
rect 14656 23962 14712 23964
rect 14736 23962 14792 23964
rect 14816 23962 14872 23964
rect 14896 23962 14952 23964
rect 14976 23962 15032 23964
rect 14656 23910 14658 23962
rect 14658 23910 14710 23962
rect 14710 23910 14712 23962
rect 14736 23910 14774 23962
rect 14774 23910 14786 23962
rect 14786 23910 14792 23962
rect 14816 23910 14838 23962
rect 14838 23910 14850 23962
rect 14850 23910 14872 23962
rect 14896 23910 14902 23962
rect 14902 23910 14914 23962
rect 14914 23910 14952 23962
rect 14976 23910 14978 23962
rect 14978 23910 15030 23962
rect 15030 23910 15032 23962
rect 14656 23908 14712 23910
rect 14736 23908 14792 23910
rect 14816 23908 14872 23910
rect 14896 23908 14952 23910
rect 14976 23908 15032 23910
rect 14656 22874 14712 22876
rect 14736 22874 14792 22876
rect 14816 22874 14872 22876
rect 14896 22874 14952 22876
rect 14976 22874 15032 22876
rect 14656 22822 14658 22874
rect 14658 22822 14710 22874
rect 14710 22822 14712 22874
rect 14736 22822 14774 22874
rect 14774 22822 14786 22874
rect 14786 22822 14792 22874
rect 14816 22822 14838 22874
rect 14838 22822 14850 22874
rect 14850 22822 14872 22874
rect 14896 22822 14902 22874
rect 14902 22822 14914 22874
rect 14914 22822 14952 22874
rect 14976 22822 14978 22874
rect 14978 22822 15030 22874
rect 15030 22822 15032 22874
rect 14656 22820 14712 22822
rect 14736 22820 14792 22822
rect 14816 22820 14872 22822
rect 14896 22820 14952 22822
rect 14976 22820 15032 22822
rect 20656 23962 20712 23964
rect 20736 23962 20792 23964
rect 20816 23962 20872 23964
rect 20896 23962 20952 23964
rect 20976 23962 21032 23964
rect 20656 23910 20658 23962
rect 20658 23910 20710 23962
rect 20710 23910 20712 23962
rect 20736 23910 20774 23962
rect 20774 23910 20786 23962
rect 20786 23910 20792 23962
rect 20816 23910 20838 23962
rect 20838 23910 20850 23962
rect 20850 23910 20872 23962
rect 20896 23910 20902 23962
rect 20902 23910 20914 23962
rect 20914 23910 20952 23962
rect 20976 23910 20978 23962
rect 20978 23910 21030 23962
rect 21030 23910 21032 23962
rect 20656 23908 20712 23910
rect 20736 23908 20792 23910
rect 20816 23908 20872 23910
rect 20896 23908 20952 23910
rect 20976 23908 21032 23910
rect 19916 23418 19972 23420
rect 19996 23418 20052 23420
rect 20076 23418 20132 23420
rect 20156 23418 20212 23420
rect 20236 23418 20292 23420
rect 19916 23366 19918 23418
rect 19918 23366 19970 23418
rect 19970 23366 19972 23418
rect 19996 23366 20034 23418
rect 20034 23366 20046 23418
rect 20046 23366 20052 23418
rect 20076 23366 20098 23418
rect 20098 23366 20110 23418
rect 20110 23366 20132 23418
rect 20156 23366 20162 23418
rect 20162 23366 20174 23418
rect 20174 23366 20212 23418
rect 20236 23366 20238 23418
rect 20238 23366 20290 23418
rect 20290 23366 20292 23418
rect 19916 23364 19972 23366
rect 19996 23364 20052 23366
rect 20076 23364 20132 23366
rect 20156 23364 20212 23366
rect 20236 23364 20292 23366
rect 20656 22874 20712 22876
rect 20736 22874 20792 22876
rect 20816 22874 20872 22876
rect 20896 22874 20952 22876
rect 20976 22874 21032 22876
rect 20656 22822 20658 22874
rect 20658 22822 20710 22874
rect 20710 22822 20712 22874
rect 20736 22822 20774 22874
rect 20774 22822 20786 22874
rect 20786 22822 20792 22874
rect 20816 22822 20838 22874
rect 20838 22822 20850 22874
rect 20850 22822 20872 22874
rect 20896 22822 20902 22874
rect 20902 22822 20914 22874
rect 20914 22822 20952 22874
rect 20976 22822 20978 22874
rect 20978 22822 21030 22874
rect 21030 22822 21032 22874
rect 20656 22820 20712 22822
rect 20736 22820 20792 22822
rect 20816 22820 20872 22822
rect 20896 22820 20952 22822
rect 20976 22820 21032 22822
rect 14656 21786 14712 21788
rect 14736 21786 14792 21788
rect 14816 21786 14872 21788
rect 14896 21786 14952 21788
rect 14976 21786 15032 21788
rect 14656 21734 14658 21786
rect 14658 21734 14710 21786
rect 14710 21734 14712 21786
rect 14736 21734 14774 21786
rect 14774 21734 14786 21786
rect 14786 21734 14792 21786
rect 14816 21734 14838 21786
rect 14838 21734 14850 21786
rect 14850 21734 14872 21786
rect 14896 21734 14902 21786
rect 14902 21734 14914 21786
rect 14914 21734 14952 21786
rect 14976 21734 14978 21786
rect 14978 21734 15030 21786
rect 15030 21734 15032 21786
rect 14656 21732 14712 21734
rect 14736 21732 14792 21734
rect 14816 21732 14872 21734
rect 14896 21732 14952 21734
rect 14976 21732 15032 21734
rect 14656 20698 14712 20700
rect 14736 20698 14792 20700
rect 14816 20698 14872 20700
rect 14896 20698 14952 20700
rect 14976 20698 15032 20700
rect 14656 20646 14658 20698
rect 14658 20646 14710 20698
rect 14710 20646 14712 20698
rect 14736 20646 14774 20698
rect 14774 20646 14786 20698
rect 14786 20646 14792 20698
rect 14816 20646 14838 20698
rect 14838 20646 14850 20698
rect 14850 20646 14872 20698
rect 14896 20646 14902 20698
rect 14902 20646 14914 20698
rect 14914 20646 14952 20698
rect 14976 20646 14978 20698
rect 14978 20646 15030 20698
rect 15030 20646 15032 20698
rect 14656 20644 14712 20646
rect 14736 20644 14792 20646
rect 14816 20644 14872 20646
rect 14896 20644 14952 20646
rect 14976 20644 15032 20646
rect 11610 13368 11666 13424
rect 11242 9560 11298 9616
rect 11242 6704 11298 6760
rect 13916 19066 13972 19068
rect 13996 19066 14052 19068
rect 14076 19066 14132 19068
rect 14156 19066 14212 19068
rect 14236 19066 14292 19068
rect 13916 19014 13918 19066
rect 13918 19014 13970 19066
rect 13970 19014 13972 19066
rect 13996 19014 14034 19066
rect 14034 19014 14046 19066
rect 14046 19014 14052 19066
rect 14076 19014 14098 19066
rect 14098 19014 14110 19066
rect 14110 19014 14132 19066
rect 14156 19014 14162 19066
rect 14162 19014 14174 19066
rect 14174 19014 14212 19066
rect 14236 19014 14238 19066
rect 14238 19014 14290 19066
rect 14290 19014 14292 19066
rect 13916 19012 13972 19014
rect 13996 19012 14052 19014
rect 14076 19012 14132 19014
rect 14156 19012 14212 19014
rect 14236 19012 14292 19014
rect 14656 19610 14712 19612
rect 14736 19610 14792 19612
rect 14816 19610 14872 19612
rect 14896 19610 14952 19612
rect 14976 19610 15032 19612
rect 14656 19558 14658 19610
rect 14658 19558 14710 19610
rect 14710 19558 14712 19610
rect 14736 19558 14774 19610
rect 14774 19558 14786 19610
rect 14786 19558 14792 19610
rect 14816 19558 14838 19610
rect 14838 19558 14850 19610
rect 14850 19558 14872 19610
rect 14896 19558 14902 19610
rect 14902 19558 14914 19610
rect 14914 19558 14952 19610
rect 14976 19558 14978 19610
rect 14978 19558 15030 19610
rect 15030 19558 15032 19610
rect 14656 19556 14712 19558
rect 14736 19556 14792 19558
rect 14816 19556 14872 19558
rect 14896 19556 14952 19558
rect 14976 19556 15032 19558
rect 14922 19352 14978 19408
rect 13916 17978 13972 17980
rect 13996 17978 14052 17980
rect 14076 17978 14132 17980
rect 14156 17978 14212 17980
rect 14236 17978 14292 17980
rect 13916 17926 13918 17978
rect 13918 17926 13970 17978
rect 13970 17926 13972 17978
rect 13996 17926 14034 17978
rect 14034 17926 14046 17978
rect 14046 17926 14052 17978
rect 14076 17926 14098 17978
rect 14098 17926 14110 17978
rect 14110 17926 14132 17978
rect 14156 17926 14162 17978
rect 14162 17926 14174 17978
rect 14174 17926 14212 17978
rect 14236 17926 14238 17978
rect 14238 17926 14290 17978
rect 14290 17926 14292 17978
rect 13916 17924 13972 17926
rect 13996 17924 14052 17926
rect 14076 17924 14132 17926
rect 14156 17924 14212 17926
rect 14236 17924 14292 17926
rect 13916 16890 13972 16892
rect 13996 16890 14052 16892
rect 14076 16890 14132 16892
rect 14156 16890 14212 16892
rect 14236 16890 14292 16892
rect 13916 16838 13918 16890
rect 13918 16838 13970 16890
rect 13970 16838 13972 16890
rect 13996 16838 14034 16890
rect 14034 16838 14046 16890
rect 14046 16838 14052 16890
rect 14076 16838 14098 16890
rect 14098 16838 14110 16890
rect 14110 16838 14132 16890
rect 14156 16838 14162 16890
rect 14162 16838 14174 16890
rect 14174 16838 14212 16890
rect 14236 16838 14238 16890
rect 14238 16838 14290 16890
rect 14290 16838 14292 16890
rect 13916 16836 13972 16838
rect 13996 16836 14052 16838
rect 14076 16836 14132 16838
rect 14156 16836 14212 16838
rect 14236 16836 14292 16838
rect 13916 15802 13972 15804
rect 13996 15802 14052 15804
rect 14076 15802 14132 15804
rect 14156 15802 14212 15804
rect 14236 15802 14292 15804
rect 13916 15750 13918 15802
rect 13918 15750 13970 15802
rect 13970 15750 13972 15802
rect 13996 15750 14034 15802
rect 14034 15750 14046 15802
rect 14046 15750 14052 15802
rect 14076 15750 14098 15802
rect 14098 15750 14110 15802
rect 14110 15750 14132 15802
rect 14156 15750 14162 15802
rect 14162 15750 14174 15802
rect 14174 15750 14212 15802
rect 14236 15750 14238 15802
rect 14238 15750 14290 15802
rect 14290 15750 14292 15802
rect 13916 15748 13972 15750
rect 13996 15748 14052 15750
rect 14076 15748 14132 15750
rect 14156 15748 14212 15750
rect 14236 15748 14292 15750
rect 13916 14714 13972 14716
rect 13996 14714 14052 14716
rect 14076 14714 14132 14716
rect 14156 14714 14212 14716
rect 14236 14714 14292 14716
rect 13916 14662 13918 14714
rect 13918 14662 13970 14714
rect 13970 14662 13972 14714
rect 13996 14662 14034 14714
rect 14034 14662 14046 14714
rect 14046 14662 14052 14714
rect 14076 14662 14098 14714
rect 14098 14662 14110 14714
rect 14110 14662 14132 14714
rect 14156 14662 14162 14714
rect 14162 14662 14174 14714
rect 14174 14662 14212 14714
rect 14236 14662 14238 14714
rect 14238 14662 14290 14714
rect 14290 14662 14292 14714
rect 13916 14660 13972 14662
rect 13996 14660 14052 14662
rect 14076 14660 14132 14662
rect 14156 14660 14212 14662
rect 14236 14660 14292 14662
rect 13916 13626 13972 13628
rect 13996 13626 14052 13628
rect 14076 13626 14132 13628
rect 14156 13626 14212 13628
rect 14236 13626 14292 13628
rect 13916 13574 13918 13626
rect 13918 13574 13970 13626
rect 13970 13574 13972 13626
rect 13996 13574 14034 13626
rect 14034 13574 14046 13626
rect 14046 13574 14052 13626
rect 14076 13574 14098 13626
rect 14098 13574 14110 13626
rect 14110 13574 14132 13626
rect 14156 13574 14162 13626
rect 14162 13574 14174 13626
rect 14174 13574 14212 13626
rect 14236 13574 14238 13626
rect 14238 13574 14290 13626
rect 14290 13574 14292 13626
rect 13916 13572 13972 13574
rect 13996 13572 14052 13574
rect 14076 13572 14132 13574
rect 14156 13572 14212 13574
rect 14236 13572 14292 13574
rect 14370 13368 14426 13424
rect 14278 12708 14334 12744
rect 14278 12688 14280 12708
rect 14280 12688 14332 12708
rect 14332 12688 14334 12708
rect 13916 12538 13972 12540
rect 13996 12538 14052 12540
rect 14076 12538 14132 12540
rect 14156 12538 14212 12540
rect 14236 12538 14292 12540
rect 13916 12486 13918 12538
rect 13918 12486 13970 12538
rect 13970 12486 13972 12538
rect 13996 12486 14034 12538
rect 14034 12486 14046 12538
rect 14046 12486 14052 12538
rect 14076 12486 14098 12538
rect 14098 12486 14110 12538
rect 14110 12486 14132 12538
rect 14156 12486 14162 12538
rect 14162 12486 14174 12538
rect 14174 12486 14212 12538
rect 14236 12486 14238 12538
rect 14238 12486 14290 12538
rect 14290 12486 14292 12538
rect 13916 12484 13972 12486
rect 13996 12484 14052 12486
rect 14076 12484 14132 12486
rect 14156 12484 14212 12486
rect 14236 12484 14292 12486
rect 13916 11450 13972 11452
rect 13996 11450 14052 11452
rect 14076 11450 14132 11452
rect 14156 11450 14212 11452
rect 14236 11450 14292 11452
rect 13916 11398 13918 11450
rect 13918 11398 13970 11450
rect 13970 11398 13972 11450
rect 13996 11398 14034 11450
rect 14034 11398 14046 11450
rect 14046 11398 14052 11450
rect 14076 11398 14098 11450
rect 14098 11398 14110 11450
rect 14110 11398 14132 11450
rect 14156 11398 14162 11450
rect 14162 11398 14174 11450
rect 14174 11398 14212 11450
rect 14236 11398 14238 11450
rect 14238 11398 14290 11450
rect 14290 11398 14292 11450
rect 13916 11396 13972 11398
rect 13996 11396 14052 11398
rect 14076 11396 14132 11398
rect 14156 11396 14212 11398
rect 14236 11396 14292 11398
rect 12622 9988 12678 10024
rect 12622 9968 12624 9988
rect 12624 9968 12676 9988
rect 12676 9968 12678 9988
rect 11886 9560 11942 9616
rect 8656 3290 8712 3292
rect 8736 3290 8792 3292
rect 8816 3290 8872 3292
rect 8896 3290 8952 3292
rect 8976 3290 9032 3292
rect 8656 3238 8658 3290
rect 8658 3238 8710 3290
rect 8710 3238 8712 3290
rect 8736 3238 8774 3290
rect 8774 3238 8786 3290
rect 8786 3238 8792 3290
rect 8816 3238 8838 3290
rect 8838 3238 8850 3290
rect 8850 3238 8872 3290
rect 8896 3238 8902 3290
rect 8902 3238 8914 3290
rect 8914 3238 8952 3290
rect 8976 3238 8978 3290
rect 8978 3238 9030 3290
rect 9030 3238 9032 3290
rect 8656 3236 8712 3238
rect 8736 3236 8792 3238
rect 8816 3236 8872 3238
rect 8896 3236 8952 3238
rect 8976 3236 9032 3238
rect 7916 2746 7972 2748
rect 7996 2746 8052 2748
rect 8076 2746 8132 2748
rect 8156 2746 8212 2748
rect 8236 2746 8292 2748
rect 7916 2694 7918 2746
rect 7918 2694 7970 2746
rect 7970 2694 7972 2746
rect 7996 2694 8034 2746
rect 8034 2694 8046 2746
rect 8046 2694 8052 2746
rect 8076 2694 8098 2746
rect 8098 2694 8110 2746
rect 8110 2694 8132 2746
rect 8156 2694 8162 2746
rect 8162 2694 8174 2746
rect 8174 2694 8212 2746
rect 8236 2694 8238 2746
rect 8238 2694 8290 2746
rect 8290 2694 8292 2746
rect 7916 2692 7972 2694
rect 7996 2692 8052 2694
rect 8076 2692 8132 2694
rect 8156 2692 8212 2694
rect 8236 2692 8292 2694
rect 2656 2202 2712 2204
rect 2736 2202 2792 2204
rect 2816 2202 2872 2204
rect 2896 2202 2952 2204
rect 2976 2202 3032 2204
rect 2656 2150 2658 2202
rect 2658 2150 2710 2202
rect 2710 2150 2712 2202
rect 2736 2150 2774 2202
rect 2774 2150 2786 2202
rect 2786 2150 2792 2202
rect 2816 2150 2838 2202
rect 2838 2150 2850 2202
rect 2850 2150 2872 2202
rect 2896 2150 2902 2202
rect 2902 2150 2914 2202
rect 2914 2150 2952 2202
rect 2976 2150 2978 2202
rect 2978 2150 3030 2202
rect 3030 2150 3032 2202
rect 2656 2148 2712 2150
rect 2736 2148 2792 2150
rect 2816 2148 2872 2150
rect 2896 2148 2952 2150
rect 2976 2148 3032 2150
rect 8656 2202 8712 2204
rect 8736 2202 8792 2204
rect 8816 2202 8872 2204
rect 8896 2202 8952 2204
rect 8976 2202 9032 2204
rect 8656 2150 8658 2202
rect 8658 2150 8710 2202
rect 8710 2150 8712 2202
rect 8736 2150 8774 2202
rect 8774 2150 8786 2202
rect 8786 2150 8792 2202
rect 8816 2150 8838 2202
rect 8838 2150 8850 2202
rect 8850 2150 8872 2202
rect 8896 2150 8902 2202
rect 8902 2150 8914 2202
rect 8914 2150 8952 2202
rect 8976 2150 8978 2202
rect 8978 2150 9030 2202
rect 9030 2150 9032 2202
rect 8656 2148 8712 2150
rect 8736 2148 8792 2150
rect 8816 2148 8872 2150
rect 8896 2148 8952 2150
rect 8976 2148 9032 2150
rect 12438 9424 12494 9480
rect 12162 7928 12218 7984
rect 14656 18522 14712 18524
rect 14736 18522 14792 18524
rect 14816 18522 14872 18524
rect 14896 18522 14952 18524
rect 14976 18522 15032 18524
rect 14656 18470 14658 18522
rect 14658 18470 14710 18522
rect 14710 18470 14712 18522
rect 14736 18470 14774 18522
rect 14774 18470 14786 18522
rect 14786 18470 14792 18522
rect 14816 18470 14838 18522
rect 14838 18470 14850 18522
rect 14850 18470 14872 18522
rect 14896 18470 14902 18522
rect 14902 18470 14914 18522
rect 14914 18470 14952 18522
rect 14976 18470 14978 18522
rect 14978 18470 15030 18522
rect 15030 18470 15032 18522
rect 14656 18468 14712 18470
rect 14736 18468 14792 18470
rect 14816 18468 14872 18470
rect 14896 18468 14952 18470
rect 14976 18468 15032 18470
rect 14656 17434 14712 17436
rect 14736 17434 14792 17436
rect 14816 17434 14872 17436
rect 14896 17434 14952 17436
rect 14976 17434 15032 17436
rect 14656 17382 14658 17434
rect 14658 17382 14710 17434
rect 14710 17382 14712 17434
rect 14736 17382 14774 17434
rect 14774 17382 14786 17434
rect 14786 17382 14792 17434
rect 14816 17382 14838 17434
rect 14838 17382 14850 17434
rect 14850 17382 14872 17434
rect 14896 17382 14902 17434
rect 14902 17382 14914 17434
rect 14914 17382 14952 17434
rect 14976 17382 14978 17434
rect 14978 17382 15030 17434
rect 15030 17382 15032 17434
rect 14656 17380 14712 17382
rect 14736 17380 14792 17382
rect 14816 17380 14872 17382
rect 14896 17380 14952 17382
rect 14976 17380 15032 17382
rect 15566 19352 15622 19408
rect 19916 22330 19972 22332
rect 19996 22330 20052 22332
rect 20076 22330 20132 22332
rect 20156 22330 20212 22332
rect 20236 22330 20292 22332
rect 19916 22278 19918 22330
rect 19918 22278 19970 22330
rect 19970 22278 19972 22330
rect 19996 22278 20034 22330
rect 20034 22278 20046 22330
rect 20046 22278 20052 22330
rect 20076 22278 20098 22330
rect 20098 22278 20110 22330
rect 20110 22278 20132 22330
rect 20156 22278 20162 22330
rect 20162 22278 20174 22330
rect 20174 22278 20212 22330
rect 20236 22278 20238 22330
rect 20238 22278 20290 22330
rect 20290 22278 20292 22330
rect 19916 22276 19972 22278
rect 19996 22276 20052 22278
rect 20076 22276 20132 22278
rect 20156 22276 20212 22278
rect 20236 22276 20292 22278
rect 20656 21786 20712 21788
rect 20736 21786 20792 21788
rect 20816 21786 20872 21788
rect 20896 21786 20952 21788
rect 20976 21786 21032 21788
rect 20656 21734 20658 21786
rect 20658 21734 20710 21786
rect 20710 21734 20712 21786
rect 20736 21734 20774 21786
rect 20774 21734 20786 21786
rect 20786 21734 20792 21786
rect 20816 21734 20838 21786
rect 20838 21734 20850 21786
rect 20850 21734 20872 21786
rect 20896 21734 20902 21786
rect 20902 21734 20914 21786
rect 20914 21734 20952 21786
rect 20976 21734 20978 21786
rect 20978 21734 21030 21786
rect 21030 21734 21032 21786
rect 20656 21732 20712 21734
rect 20736 21732 20792 21734
rect 20816 21732 20872 21734
rect 20896 21732 20952 21734
rect 20976 21732 21032 21734
rect 14656 16346 14712 16348
rect 14736 16346 14792 16348
rect 14816 16346 14872 16348
rect 14896 16346 14952 16348
rect 14976 16346 15032 16348
rect 14656 16294 14658 16346
rect 14658 16294 14710 16346
rect 14710 16294 14712 16346
rect 14736 16294 14774 16346
rect 14774 16294 14786 16346
rect 14786 16294 14792 16346
rect 14816 16294 14838 16346
rect 14838 16294 14850 16346
rect 14850 16294 14872 16346
rect 14896 16294 14902 16346
rect 14902 16294 14914 16346
rect 14914 16294 14952 16346
rect 14976 16294 14978 16346
rect 14978 16294 15030 16346
rect 15030 16294 15032 16346
rect 14656 16292 14712 16294
rect 14736 16292 14792 16294
rect 14816 16292 14872 16294
rect 14896 16292 14952 16294
rect 14976 16292 15032 16294
rect 14656 15258 14712 15260
rect 14736 15258 14792 15260
rect 14816 15258 14872 15260
rect 14896 15258 14952 15260
rect 14976 15258 15032 15260
rect 14656 15206 14658 15258
rect 14658 15206 14710 15258
rect 14710 15206 14712 15258
rect 14736 15206 14774 15258
rect 14774 15206 14786 15258
rect 14786 15206 14792 15258
rect 14816 15206 14838 15258
rect 14838 15206 14850 15258
rect 14850 15206 14872 15258
rect 14896 15206 14902 15258
rect 14902 15206 14914 15258
rect 14914 15206 14952 15258
rect 14976 15206 14978 15258
rect 14978 15206 15030 15258
rect 15030 15206 15032 15258
rect 14656 15204 14712 15206
rect 14736 15204 14792 15206
rect 14816 15204 14872 15206
rect 14896 15204 14952 15206
rect 14976 15204 15032 15206
rect 14656 14170 14712 14172
rect 14736 14170 14792 14172
rect 14816 14170 14872 14172
rect 14896 14170 14952 14172
rect 14976 14170 15032 14172
rect 14656 14118 14658 14170
rect 14658 14118 14710 14170
rect 14710 14118 14712 14170
rect 14736 14118 14774 14170
rect 14774 14118 14786 14170
rect 14786 14118 14792 14170
rect 14816 14118 14838 14170
rect 14838 14118 14850 14170
rect 14850 14118 14872 14170
rect 14896 14118 14902 14170
rect 14902 14118 14914 14170
rect 14914 14118 14952 14170
rect 14976 14118 14978 14170
rect 14978 14118 15030 14170
rect 15030 14118 15032 14170
rect 14656 14116 14712 14118
rect 14736 14116 14792 14118
rect 14816 14116 14872 14118
rect 14896 14116 14952 14118
rect 14976 14116 15032 14118
rect 14656 13082 14712 13084
rect 14736 13082 14792 13084
rect 14816 13082 14872 13084
rect 14896 13082 14952 13084
rect 14976 13082 15032 13084
rect 14656 13030 14658 13082
rect 14658 13030 14710 13082
rect 14710 13030 14712 13082
rect 14736 13030 14774 13082
rect 14774 13030 14786 13082
rect 14786 13030 14792 13082
rect 14816 13030 14838 13082
rect 14838 13030 14850 13082
rect 14850 13030 14872 13082
rect 14896 13030 14902 13082
rect 14902 13030 14914 13082
rect 14914 13030 14952 13082
rect 14976 13030 14978 13082
rect 14978 13030 15030 13082
rect 15030 13030 15032 13082
rect 14656 13028 14712 13030
rect 14736 13028 14792 13030
rect 14816 13028 14872 13030
rect 14896 13028 14952 13030
rect 14976 13028 15032 13030
rect 14656 11994 14712 11996
rect 14736 11994 14792 11996
rect 14816 11994 14872 11996
rect 14896 11994 14952 11996
rect 14976 11994 15032 11996
rect 14656 11942 14658 11994
rect 14658 11942 14710 11994
rect 14710 11942 14712 11994
rect 14736 11942 14774 11994
rect 14774 11942 14786 11994
rect 14786 11942 14792 11994
rect 14816 11942 14838 11994
rect 14838 11942 14850 11994
rect 14850 11942 14872 11994
rect 14896 11942 14902 11994
rect 14902 11942 14914 11994
rect 14914 11942 14952 11994
rect 14976 11942 14978 11994
rect 14978 11942 15030 11994
rect 15030 11942 15032 11994
rect 14656 11940 14712 11942
rect 14736 11940 14792 11942
rect 14816 11940 14872 11942
rect 14896 11940 14952 11942
rect 14976 11940 15032 11942
rect 14462 11600 14518 11656
rect 14656 10906 14712 10908
rect 14736 10906 14792 10908
rect 14816 10906 14872 10908
rect 14896 10906 14952 10908
rect 14976 10906 15032 10908
rect 14656 10854 14658 10906
rect 14658 10854 14710 10906
rect 14710 10854 14712 10906
rect 14736 10854 14774 10906
rect 14774 10854 14786 10906
rect 14786 10854 14792 10906
rect 14816 10854 14838 10906
rect 14838 10854 14850 10906
rect 14850 10854 14872 10906
rect 14896 10854 14902 10906
rect 14902 10854 14914 10906
rect 14914 10854 14952 10906
rect 14976 10854 14978 10906
rect 14978 10854 15030 10906
rect 15030 10854 15032 10906
rect 14656 10852 14712 10854
rect 14736 10852 14792 10854
rect 14816 10852 14872 10854
rect 14896 10852 14952 10854
rect 14976 10852 15032 10854
rect 13916 10362 13972 10364
rect 13996 10362 14052 10364
rect 14076 10362 14132 10364
rect 14156 10362 14212 10364
rect 14236 10362 14292 10364
rect 13916 10310 13918 10362
rect 13918 10310 13970 10362
rect 13970 10310 13972 10362
rect 13996 10310 14034 10362
rect 14034 10310 14046 10362
rect 14046 10310 14052 10362
rect 14076 10310 14098 10362
rect 14098 10310 14110 10362
rect 14110 10310 14132 10362
rect 14156 10310 14162 10362
rect 14162 10310 14174 10362
rect 14174 10310 14212 10362
rect 14236 10310 14238 10362
rect 14238 10310 14290 10362
rect 14290 10310 14292 10362
rect 13916 10308 13972 10310
rect 13996 10308 14052 10310
rect 14076 10308 14132 10310
rect 14156 10308 14212 10310
rect 14236 10308 14292 10310
rect 13916 9274 13972 9276
rect 13996 9274 14052 9276
rect 14076 9274 14132 9276
rect 14156 9274 14212 9276
rect 14236 9274 14292 9276
rect 13916 9222 13918 9274
rect 13918 9222 13970 9274
rect 13970 9222 13972 9274
rect 13996 9222 14034 9274
rect 14034 9222 14046 9274
rect 14046 9222 14052 9274
rect 14076 9222 14098 9274
rect 14098 9222 14110 9274
rect 14110 9222 14132 9274
rect 14156 9222 14162 9274
rect 14162 9222 14174 9274
rect 14174 9222 14212 9274
rect 14236 9222 14238 9274
rect 14238 9222 14290 9274
rect 14290 9222 14292 9274
rect 13916 9220 13972 9222
rect 13996 9220 14052 9222
rect 14076 9220 14132 9222
rect 14156 9220 14212 9222
rect 14236 9220 14292 9222
rect 13916 8186 13972 8188
rect 13996 8186 14052 8188
rect 14076 8186 14132 8188
rect 14156 8186 14212 8188
rect 14236 8186 14292 8188
rect 13916 8134 13918 8186
rect 13918 8134 13970 8186
rect 13970 8134 13972 8186
rect 13996 8134 14034 8186
rect 14034 8134 14046 8186
rect 14046 8134 14052 8186
rect 14076 8134 14098 8186
rect 14098 8134 14110 8186
rect 14110 8134 14132 8186
rect 14156 8134 14162 8186
rect 14162 8134 14174 8186
rect 14174 8134 14212 8186
rect 14236 8134 14238 8186
rect 14238 8134 14290 8186
rect 14290 8134 14292 8186
rect 13916 8132 13972 8134
rect 13996 8132 14052 8134
rect 14076 8132 14132 8134
rect 14156 8132 14212 8134
rect 14236 8132 14292 8134
rect 14656 9818 14712 9820
rect 14736 9818 14792 9820
rect 14816 9818 14872 9820
rect 14896 9818 14952 9820
rect 14976 9818 15032 9820
rect 14656 9766 14658 9818
rect 14658 9766 14710 9818
rect 14710 9766 14712 9818
rect 14736 9766 14774 9818
rect 14774 9766 14786 9818
rect 14786 9766 14792 9818
rect 14816 9766 14838 9818
rect 14838 9766 14850 9818
rect 14850 9766 14872 9818
rect 14896 9766 14902 9818
rect 14902 9766 14914 9818
rect 14914 9766 14952 9818
rect 14976 9766 14978 9818
rect 14978 9766 15030 9818
rect 15030 9766 15032 9818
rect 14656 9764 14712 9766
rect 14736 9764 14792 9766
rect 14816 9764 14872 9766
rect 14896 9764 14952 9766
rect 14976 9764 15032 9766
rect 13916 7098 13972 7100
rect 13996 7098 14052 7100
rect 14076 7098 14132 7100
rect 14156 7098 14212 7100
rect 14236 7098 14292 7100
rect 13916 7046 13918 7098
rect 13918 7046 13970 7098
rect 13970 7046 13972 7098
rect 13996 7046 14034 7098
rect 14034 7046 14046 7098
rect 14046 7046 14052 7098
rect 14076 7046 14098 7098
rect 14098 7046 14110 7098
rect 14110 7046 14132 7098
rect 14156 7046 14162 7098
rect 14162 7046 14174 7098
rect 14174 7046 14212 7098
rect 14236 7046 14238 7098
rect 14238 7046 14290 7098
rect 14290 7046 14292 7098
rect 13916 7044 13972 7046
rect 13996 7044 14052 7046
rect 14076 7044 14132 7046
rect 14156 7044 14212 7046
rect 14236 7044 14292 7046
rect 13916 6010 13972 6012
rect 13996 6010 14052 6012
rect 14076 6010 14132 6012
rect 14156 6010 14212 6012
rect 14236 6010 14292 6012
rect 13916 5958 13918 6010
rect 13918 5958 13970 6010
rect 13970 5958 13972 6010
rect 13996 5958 14034 6010
rect 14034 5958 14046 6010
rect 14046 5958 14052 6010
rect 14076 5958 14098 6010
rect 14098 5958 14110 6010
rect 14110 5958 14132 6010
rect 14156 5958 14162 6010
rect 14162 5958 14174 6010
rect 14174 5958 14212 6010
rect 14236 5958 14238 6010
rect 14238 5958 14290 6010
rect 14290 5958 14292 6010
rect 13916 5956 13972 5958
rect 13996 5956 14052 5958
rect 14076 5956 14132 5958
rect 14156 5956 14212 5958
rect 14236 5956 14292 5958
rect 13916 4922 13972 4924
rect 13996 4922 14052 4924
rect 14076 4922 14132 4924
rect 14156 4922 14212 4924
rect 14236 4922 14292 4924
rect 13916 4870 13918 4922
rect 13918 4870 13970 4922
rect 13970 4870 13972 4922
rect 13996 4870 14034 4922
rect 14034 4870 14046 4922
rect 14046 4870 14052 4922
rect 14076 4870 14098 4922
rect 14098 4870 14110 4922
rect 14110 4870 14132 4922
rect 14156 4870 14162 4922
rect 14162 4870 14174 4922
rect 14174 4870 14212 4922
rect 14236 4870 14238 4922
rect 14238 4870 14290 4922
rect 14290 4870 14292 4922
rect 13916 4868 13972 4870
rect 13996 4868 14052 4870
rect 14076 4868 14132 4870
rect 14156 4868 14212 4870
rect 14236 4868 14292 4870
rect 14656 8730 14712 8732
rect 14736 8730 14792 8732
rect 14816 8730 14872 8732
rect 14896 8730 14952 8732
rect 14976 8730 15032 8732
rect 14656 8678 14658 8730
rect 14658 8678 14710 8730
rect 14710 8678 14712 8730
rect 14736 8678 14774 8730
rect 14774 8678 14786 8730
rect 14786 8678 14792 8730
rect 14816 8678 14838 8730
rect 14838 8678 14850 8730
rect 14850 8678 14872 8730
rect 14896 8678 14902 8730
rect 14902 8678 14914 8730
rect 14914 8678 14952 8730
rect 14976 8678 14978 8730
rect 14978 8678 15030 8730
rect 15030 8678 15032 8730
rect 14656 8676 14712 8678
rect 14736 8676 14792 8678
rect 14816 8676 14872 8678
rect 14896 8676 14952 8678
rect 14976 8676 15032 8678
rect 19916 21242 19972 21244
rect 19996 21242 20052 21244
rect 20076 21242 20132 21244
rect 20156 21242 20212 21244
rect 20236 21242 20292 21244
rect 19916 21190 19918 21242
rect 19918 21190 19970 21242
rect 19970 21190 19972 21242
rect 19996 21190 20034 21242
rect 20034 21190 20046 21242
rect 20046 21190 20052 21242
rect 20076 21190 20098 21242
rect 20098 21190 20110 21242
rect 20110 21190 20132 21242
rect 20156 21190 20162 21242
rect 20162 21190 20174 21242
rect 20174 21190 20212 21242
rect 20236 21190 20238 21242
rect 20238 21190 20290 21242
rect 20290 21190 20292 21242
rect 19916 21188 19972 21190
rect 19996 21188 20052 21190
rect 20076 21188 20132 21190
rect 20156 21188 20212 21190
rect 20236 21188 20292 21190
rect 20656 20698 20712 20700
rect 20736 20698 20792 20700
rect 20816 20698 20872 20700
rect 20896 20698 20952 20700
rect 20976 20698 21032 20700
rect 20656 20646 20658 20698
rect 20658 20646 20710 20698
rect 20710 20646 20712 20698
rect 20736 20646 20774 20698
rect 20774 20646 20786 20698
rect 20786 20646 20792 20698
rect 20816 20646 20838 20698
rect 20838 20646 20850 20698
rect 20850 20646 20872 20698
rect 20896 20646 20902 20698
rect 20902 20646 20914 20698
rect 20914 20646 20952 20698
rect 20976 20646 20978 20698
rect 20978 20646 21030 20698
rect 21030 20646 21032 20698
rect 20656 20644 20712 20646
rect 20736 20644 20792 20646
rect 20816 20644 20872 20646
rect 20896 20644 20952 20646
rect 20976 20644 21032 20646
rect 15474 9968 15530 10024
rect 14656 7642 14712 7644
rect 14736 7642 14792 7644
rect 14816 7642 14872 7644
rect 14896 7642 14952 7644
rect 14976 7642 15032 7644
rect 14656 7590 14658 7642
rect 14658 7590 14710 7642
rect 14710 7590 14712 7642
rect 14736 7590 14774 7642
rect 14774 7590 14786 7642
rect 14786 7590 14792 7642
rect 14816 7590 14838 7642
rect 14838 7590 14850 7642
rect 14850 7590 14872 7642
rect 14896 7590 14902 7642
rect 14902 7590 14914 7642
rect 14914 7590 14952 7642
rect 14976 7590 14978 7642
rect 14978 7590 15030 7642
rect 15030 7590 15032 7642
rect 14656 7588 14712 7590
rect 14736 7588 14792 7590
rect 14816 7588 14872 7590
rect 14896 7588 14952 7590
rect 14976 7588 15032 7590
rect 14656 6554 14712 6556
rect 14736 6554 14792 6556
rect 14816 6554 14872 6556
rect 14896 6554 14952 6556
rect 14976 6554 15032 6556
rect 14656 6502 14658 6554
rect 14658 6502 14710 6554
rect 14710 6502 14712 6554
rect 14736 6502 14774 6554
rect 14774 6502 14786 6554
rect 14786 6502 14792 6554
rect 14816 6502 14838 6554
rect 14838 6502 14850 6554
rect 14850 6502 14872 6554
rect 14896 6502 14902 6554
rect 14902 6502 14914 6554
rect 14914 6502 14952 6554
rect 14976 6502 14978 6554
rect 14978 6502 15030 6554
rect 15030 6502 15032 6554
rect 14656 6500 14712 6502
rect 14736 6500 14792 6502
rect 14816 6500 14872 6502
rect 14896 6500 14952 6502
rect 14976 6500 15032 6502
rect 14656 5466 14712 5468
rect 14736 5466 14792 5468
rect 14816 5466 14872 5468
rect 14896 5466 14952 5468
rect 14976 5466 15032 5468
rect 14656 5414 14658 5466
rect 14658 5414 14710 5466
rect 14710 5414 14712 5466
rect 14736 5414 14774 5466
rect 14774 5414 14786 5466
rect 14786 5414 14792 5466
rect 14816 5414 14838 5466
rect 14838 5414 14850 5466
rect 14850 5414 14872 5466
rect 14896 5414 14902 5466
rect 14902 5414 14914 5466
rect 14914 5414 14952 5466
rect 14976 5414 14978 5466
rect 14978 5414 15030 5466
rect 15030 5414 15032 5466
rect 14656 5412 14712 5414
rect 14736 5412 14792 5414
rect 14816 5412 14872 5414
rect 14896 5412 14952 5414
rect 14976 5412 15032 5414
rect 17222 12688 17278 12744
rect 19916 20154 19972 20156
rect 19996 20154 20052 20156
rect 20076 20154 20132 20156
rect 20156 20154 20212 20156
rect 20236 20154 20292 20156
rect 19916 20102 19918 20154
rect 19918 20102 19970 20154
rect 19970 20102 19972 20154
rect 19996 20102 20034 20154
rect 20034 20102 20046 20154
rect 20046 20102 20052 20154
rect 20076 20102 20098 20154
rect 20098 20102 20110 20154
rect 20110 20102 20132 20154
rect 20156 20102 20162 20154
rect 20162 20102 20174 20154
rect 20174 20102 20212 20154
rect 20236 20102 20238 20154
rect 20238 20102 20290 20154
rect 20290 20102 20292 20154
rect 19916 20100 19972 20102
rect 19996 20100 20052 20102
rect 20076 20100 20132 20102
rect 20156 20100 20212 20102
rect 20236 20100 20292 20102
rect 20656 19610 20712 19612
rect 20736 19610 20792 19612
rect 20816 19610 20872 19612
rect 20896 19610 20952 19612
rect 20976 19610 21032 19612
rect 20656 19558 20658 19610
rect 20658 19558 20710 19610
rect 20710 19558 20712 19610
rect 20736 19558 20774 19610
rect 20774 19558 20786 19610
rect 20786 19558 20792 19610
rect 20816 19558 20838 19610
rect 20838 19558 20850 19610
rect 20850 19558 20872 19610
rect 20896 19558 20902 19610
rect 20902 19558 20914 19610
rect 20914 19558 20952 19610
rect 20976 19558 20978 19610
rect 20978 19558 21030 19610
rect 21030 19558 21032 19610
rect 20656 19556 20712 19558
rect 20736 19556 20792 19558
rect 20816 19556 20872 19558
rect 20896 19556 20952 19558
rect 20976 19556 21032 19558
rect 19916 19066 19972 19068
rect 19996 19066 20052 19068
rect 20076 19066 20132 19068
rect 20156 19066 20212 19068
rect 20236 19066 20292 19068
rect 19916 19014 19918 19066
rect 19918 19014 19970 19066
rect 19970 19014 19972 19066
rect 19996 19014 20034 19066
rect 20034 19014 20046 19066
rect 20046 19014 20052 19066
rect 20076 19014 20098 19066
rect 20098 19014 20110 19066
rect 20110 19014 20132 19066
rect 20156 19014 20162 19066
rect 20162 19014 20174 19066
rect 20174 19014 20212 19066
rect 20236 19014 20238 19066
rect 20238 19014 20290 19066
rect 20290 19014 20292 19066
rect 19916 19012 19972 19014
rect 19996 19012 20052 19014
rect 20076 19012 20132 19014
rect 20156 19012 20212 19014
rect 20236 19012 20292 19014
rect 23294 19080 23350 19136
rect 20656 18522 20712 18524
rect 20736 18522 20792 18524
rect 20816 18522 20872 18524
rect 20896 18522 20952 18524
rect 20976 18522 21032 18524
rect 20656 18470 20658 18522
rect 20658 18470 20710 18522
rect 20710 18470 20712 18522
rect 20736 18470 20774 18522
rect 20774 18470 20786 18522
rect 20786 18470 20792 18522
rect 20816 18470 20838 18522
rect 20838 18470 20850 18522
rect 20850 18470 20872 18522
rect 20896 18470 20902 18522
rect 20902 18470 20914 18522
rect 20914 18470 20952 18522
rect 20976 18470 20978 18522
rect 20978 18470 21030 18522
rect 21030 18470 21032 18522
rect 20656 18468 20712 18470
rect 20736 18468 20792 18470
rect 20816 18468 20872 18470
rect 20896 18468 20952 18470
rect 20976 18468 21032 18470
rect 23294 18400 23350 18456
rect 19916 17978 19972 17980
rect 19996 17978 20052 17980
rect 20076 17978 20132 17980
rect 20156 17978 20212 17980
rect 20236 17978 20292 17980
rect 19916 17926 19918 17978
rect 19918 17926 19970 17978
rect 19970 17926 19972 17978
rect 19996 17926 20034 17978
rect 20034 17926 20046 17978
rect 20046 17926 20052 17978
rect 20076 17926 20098 17978
rect 20098 17926 20110 17978
rect 20110 17926 20132 17978
rect 20156 17926 20162 17978
rect 20162 17926 20174 17978
rect 20174 17926 20212 17978
rect 20236 17926 20238 17978
rect 20238 17926 20290 17978
rect 20290 17926 20292 17978
rect 19916 17924 19972 17926
rect 19996 17924 20052 17926
rect 20076 17924 20132 17926
rect 20156 17924 20212 17926
rect 20236 17924 20292 17926
rect 20656 17434 20712 17436
rect 20736 17434 20792 17436
rect 20816 17434 20872 17436
rect 20896 17434 20952 17436
rect 20976 17434 21032 17436
rect 20656 17382 20658 17434
rect 20658 17382 20710 17434
rect 20710 17382 20712 17434
rect 20736 17382 20774 17434
rect 20774 17382 20786 17434
rect 20786 17382 20792 17434
rect 20816 17382 20838 17434
rect 20838 17382 20850 17434
rect 20850 17382 20872 17434
rect 20896 17382 20902 17434
rect 20902 17382 20914 17434
rect 20914 17382 20952 17434
rect 20976 17382 20978 17434
rect 20978 17382 21030 17434
rect 21030 17382 21032 17434
rect 20656 17380 20712 17382
rect 20736 17380 20792 17382
rect 20816 17380 20872 17382
rect 20896 17380 20952 17382
rect 20976 17380 21032 17382
rect 19916 16890 19972 16892
rect 19996 16890 20052 16892
rect 20076 16890 20132 16892
rect 20156 16890 20212 16892
rect 20236 16890 20292 16892
rect 19916 16838 19918 16890
rect 19918 16838 19970 16890
rect 19970 16838 19972 16890
rect 19996 16838 20034 16890
rect 20034 16838 20046 16890
rect 20046 16838 20052 16890
rect 20076 16838 20098 16890
rect 20098 16838 20110 16890
rect 20110 16838 20132 16890
rect 20156 16838 20162 16890
rect 20162 16838 20174 16890
rect 20174 16838 20212 16890
rect 20236 16838 20238 16890
rect 20238 16838 20290 16890
rect 20290 16838 20292 16890
rect 19916 16836 19972 16838
rect 19996 16836 20052 16838
rect 20076 16836 20132 16838
rect 20156 16836 20212 16838
rect 20236 16836 20292 16838
rect 20656 16346 20712 16348
rect 20736 16346 20792 16348
rect 20816 16346 20872 16348
rect 20896 16346 20952 16348
rect 20976 16346 21032 16348
rect 20656 16294 20658 16346
rect 20658 16294 20710 16346
rect 20710 16294 20712 16346
rect 20736 16294 20774 16346
rect 20774 16294 20786 16346
rect 20786 16294 20792 16346
rect 20816 16294 20838 16346
rect 20838 16294 20850 16346
rect 20850 16294 20872 16346
rect 20896 16294 20902 16346
rect 20902 16294 20914 16346
rect 20914 16294 20952 16346
rect 20976 16294 20978 16346
rect 20978 16294 21030 16346
rect 21030 16294 21032 16346
rect 20656 16292 20712 16294
rect 20736 16292 20792 16294
rect 20816 16292 20872 16294
rect 20896 16292 20952 16294
rect 20976 16292 21032 16294
rect 19916 15802 19972 15804
rect 19996 15802 20052 15804
rect 20076 15802 20132 15804
rect 20156 15802 20212 15804
rect 20236 15802 20292 15804
rect 19916 15750 19918 15802
rect 19918 15750 19970 15802
rect 19970 15750 19972 15802
rect 19996 15750 20034 15802
rect 20034 15750 20046 15802
rect 20046 15750 20052 15802
rect 20076 15750 20098 15802
rect 20098 15750 20110 15802
rect 20110 15750 20132 15802
rect 20156 15750 20162 15802
rect 20162 15750 20174 15802
rect 20174 15750 20212 15802
rect 20236 15750 20238 15802
rect 20238 15750 20290 15802
rect 20290 15750 20292 15802
rect 19916 15748 19972 15750
rect 19996 15748 20052 15750
rect 20076 15748 20132 15750
rect 20156 15748 20212 15750
rect 20236 15748 20292 15750
rect 19916 14714 19972 14716
rect 19996 14714 20052 14716
rect 20076 14714 20132 14716
rect 20156 14714 20212 14716
rect 20236 14714 20292 14716
rect 19916 14662 19918 14714
rect 19918 14662 19970 14714
rect 19970 14662 19972 14714
rect 19996 14662 20034 14714
rect 20034 14662 20046 14714
rect 20046 14662 20052 14714
rect 20076 14662 20098 14714
rect 20098 14662 20110 14714
rect 20110 14662 20132 14714
rect 20156 14662 20162 14714
rect 20162 14662 20174 14714
rect 20174 14662 20212 14714
rect 20236 14662 20238 14714
rect 20238 14662 20290 14714
rect 20290 14662 20292 14714
rect 19916 14660 19972 14662
rect 19996 14660 20052 14662
rect 20076 14660 20132 14662
rect 20156 14660 20212 14662
rect 20236 14660 20292 14662
rect 20656 15258 20712 15260
rect 20736 15258 20792 15260
rect 20816 15258 20872 15260
rect 20896 15258 20952 15260
rect 20976 15258 21032 15260
rect 20656 15206 20658 15258
rect 20658 15206 20710 15258
rect 20710 15206 20712 15258
rect 20736 15206 20774 15258
rect 20774 15206 20786 15258
rect 20786 15206 20792 15258
rect 20816 15206 20838 15258
rect 20838 15206 20850 15258
rect 20850 15206 20872 15258
rect 20896 15206 20902 15258
rect 20902 15206 20914 15258
rect 20914 15206 20952 15258
rect 20976 15206 20978 15258
rect 20978 15206 21030 15258
rect 21030 15206 21032 15258
rect 20656 15204 20712 15206
rect 20736 15204 20792 15206
rect 20816 15204 20872 15206
rect 20896 15204 20952 15206
rect 20976 15204 21032 15206
rect 14656 4378 14712 4380
rect 14736 4378 14792 4380
rect 14816 4378 14872 4380
rect 14896 4378 14952 4380
rect 14976 4378 15032 4380
rect 14656 4326 14658 4378
rect 14658 4326 14710 4378
rect 14710 4326 14712 4378
rect 14736 4326 14774 4378
rect 14774 4326 14786 4378
rect 14786 4326 14792 4378
rect 14816 4326 14838 4378
rect 14838 4326 14850 4378
rect 14850 4326 14872 4378
rect 14896 4326 14902 4378
rect 14902 4326 14914 4378
rect 14914 4326 14952 4378
rect 14976 4326 14978 4378
rect 14978 4326 15030 4378
rect 15030 4326 15032 4378
rect 14656 4324 14712 4326
rect 14736 4324 14792 4326
rect 14816 4324 14872 4326
rect 14896 4324 14952 4326
rect 14976 4324 15032 4326
rect 13916 3834 13972 3836
rect 13996 3834 14052 3836
rect 14076 3834 14132 3836
rect 14156 3834 14212 3836
rect 14236 3834 14292 3836
rect 13916 3782 13918 3834
rect 13918 3782 13970 3834
rect 13970 3782 13972 3834
rect 13996 3782 14034 3834
rect 14034 3782 14046 3834
rect 14046 3782 14052 3834
rect 14076 3782 14098 3834
rect 14098 3782 14110 3834
rect 14110 3782 14132 3834
rect 14156 3782 14162 3834
rect 14162 3782 14174 3834
rect 14174 3782 14212 3834
rect 14236 3782 14238 3834
rect 14238 3782 14290 3834
rect 14290 3782 14292 3834
rect 13916 3780 13972 3782
rect 13996 3780 14052 3782
rect 14076 3780 14132 3782
rect 14156 3780 14212 3782
rect 14236 3780 14292 3782
rect 14656 3290 14712 3292
rect 14736 3290 14792 3292
rect 14816 3290 14872 3292
rect 14896 3290 14952 3292
rect 14976 3290 15032 3292
rect 14656 3238 14658 3290
rect 14658 3238 14710 3290
rect 14710 3238 14712 3290
rect 14736 3238 14774 3290
rect 14774 3238 14786 3290
rect 14786 3238 14792 3290
rect 14816 3238 14838 3290
rect 14838 3238 14850 3290
rect 14850 3238 14872 3290
rect 14896 3238 14902 3290
rect 14902 3238 14914 3290
rect 14914 3238 14952 3290
rect 14976 3238 14978 3290
rect 14978 3238 15030 3290
rect 15030 3238 15032 3290
rect 14656 3236 14712 3238
rect 14736 3236 14792 3238
rect 14816 3236 14872 3238
rect 14896 3236 14952 3238
rect 14976 3236 15032 3238
rect 13916 2746 13972 2748
rect 13996 2746 14052 2748
rect 14076 2746 14132 2748
rect 14156 2746 14212 2748
rect 14236 2746 14292 2748
rect 13916 2694 13918 2746
rect 13918 2694 13970 2746
rect 13970 2694 13972 2746
rect 13996 2694 14034 2746
rect 14034 2694 14046 2746
rect 14046 2694 14052 2746
rect 14076 2694 14098 2746
rect 14098 2694 14110 2746
rect 14110 2694 14132 2746
rect 14156 2694 14162 2746
rect 14162 2694 14174 2746
rect 14174 2694 14212 2746
rect 14236 2694 14238 2746
rect 14238 2694 14290 2746
rect 14290 2694 14292 2746
rect 13916 2692 13972 2694
rect 13996 2692 14052 2694
rect 14076 2692 14132 2694
rect 14156 2692 14212 2694
rect 14236 2692 14292 2694
rect 19916 13626 19972 13628
rect 19996 13626 20052 13628
rect 20076 13626 20132 13628
rect 20156 13626 20212 13628
rect 20236 13626 20292 13628
rect 19916 13574 19918 13626
rect 19918 13574 19970 13626
rect 19970 13574 19972 13626
rect 19996 13574 20034 13626
rect 20034 13574 20046 13626
rect 20046 13574 20052 13626
rect 20076 13574 20098 13626
rect 20098 13574 20110 13626
rect 20110 13574 20132 13626
rect 20156 13574 20162 13626
rect 20162 13574 20174 13626
rect 20174 13574 20212 13626
rect 20236 13574 20238 13626
rect 20238 13574 20290 13626
rect 20290 13574 20292 13626
rect 19916 13572 19972 13574
rect 19996 13572 20052 13574
rect 20076 13572 20132 13574
rect 20156 13572 20212 13574
rect 20236 13572 20292 13574
rect 20656 14170 20712 14172
rect 20736 14170 20792 14172
rect 20816 14170 20872 14172
rect 20896 14170 20952 14172
rect 20976 14170 21032 14172
rect 20656 14118 20658 14170
rect 20658 14118 20710 14170
rect 20710 14118 20712 14170
rect 20736 14118 20774 14170
rect 20774 14118 20786 14170
rect 20786 14118 20792 14170
rect 20816 14118 20838 14170
rect 20838 14118 20850 14170
rect 20850 14118 20872 14170
rect 20896 14118 20902 14170
rect 20902 14118 20914 14170
rect 20914 14118 20952 14170
rect 20976 14118 20978 14170
rect 20978 14118 21030 14170
rect 21030 14118 21032 14170
rect 20656 14116 20712 14118
rect 20736 14116 20792 14118
rect 20816 14116 20872 14118
rect 20896 14116 20952 14118
rect 20976 14116 21032 14118
rect 20656 13082 20712 13084
rect 20736 13082 20792 13084
rect 20816 13082 20872 13084
rect 20896 13082 20952 13084
rect 20976 13082 21032 13084
rect 20656 13030 20658 13082
rect 20658 13030 20710 13082
rect 20710 13030 20712 13082
rect 20736 13030 20774 13082
rect 20774 13030 20786 13082
rect 20786 13030 20792 13082
rect 20816 13030 20838 13082
rect 20838 13030 20850 13082
rect 20850 13030 20872 13082
rect 20896 13030 20902 13082
rect 20902 13030 20914 13082
rect 20914 13030 20952 13082
rect 20976 13030 20978 13082
rect 20978 13030 21030 13082
rect 21030 13030 21032 13082
rect 20656 13028 20712 13030
rect 20736 13028 20792 13030
rect 20816 13028 20872 13030
rect 20896 13028 20952 13030
rect 20976 13028 21032 13030
rect 21546 13368 21602 13424
rect 19916 12538 19972 12540
rect 19996 12538 20052 12540
rect 20076 12538 20132 12540
rect 20156 12538 20212 12540
rect 20236 12538 20292 12540
rect 19916 12486 19918 12538
rect 19918 12486 19970 12538
rect 19970 12486 19972 12538
rect 19996 12486 20034 12538
rect 20034 12486 20046 12538
rect 20046 12486 20052 12538
rect 20076 12486 20098 12538
rect 20098 12486 20110 12538
rect 20110 12486 20132 12538
rect 20156 12486 20162 12538
rect 20162 12486 20174 12538
rect 20174 12486 20212 12538
rect 20236 12486 20238 12538
rect 20238 12486 20290 12538
rect 20290 12486 20292 12538
rect 19916 12484 19972 12486
rect 19996 12484 20052 12486
rect 20076 12484 20132 12486
rect 20156 12484 20212 12486
rect 20236 12484 20292 12486
rect 19916 11450 19972 11452
rect 19996 11450 20052 11452
rect 20076 11450 20132 11452
rect 20156 11450 20212 11452
rect 20236 11450 20292 11452
rect 19916 11398 19918 11450
rect 19918 11398 19970 11450
rect 19970 11398 19972 11450
rect 19996 11398 20034 11450
rect 20034 11398 20046 11450
rect 20046 11398 20052 11450
rect 20076 11398 20098 11450
rect 20098 11398 20110 11450
rect 20110 11398 20132 11450
rect 20156 11398 20162 11450
rect 20162 11398 20174 11450
rect 20174 11398 20212 11450
rect 20236 11398 20238 11450
rect 20238 11398 20290 11450
rect 20290 11398 20292 11450
rect 19916 11396 19972 11398
rect 19996 11396 20052 11398
rect 20076 11396 20132 11398
rect 20156 11396 20212 11398
rect 20236 11396 20292 11398
rect 19798 10512 19854 10568
rect 19916 10362 19972 10364
rect 19996 10362 20052 10364
rect 20076 10362 20132 10364
rect 20156 10362 20212 10364
rect 20236 10362 20292 10364
rect 19916 10310 19918 10362
rect 19918 10310 19970 10362
rect 19970 10310 19972 10362
rect 19996 10310 20034 10362
rect 20034 10310 20046 10362
rect 20046 10310 20052 10362
rect 20076 10310 20098 10362
rect 20098 10310 20110 10362
rect 20110 10310 20132 10362
rect 20156 10310 20162 10362
rect 20162 10310 20174 10362
rect 20174 10310 20212 10362
rect 20236 10310 20238 10362
rect 20238 10310 20290 10362
rect 20290 10310 20292 10362
rect 19916 10308 19972 10310
rect 19996 10308 20052 10310
rect 20076 10308 20132 10310
rect 20156 10308 20212 10310
rect 20236 10308 20292 10310
rect 20656 11994 20712 11996
rect 20736 11994 20792 11996
rect 20816 11994 20872 11996
rect 20896 11994 20952 11996
rect 20976 11994 21032 11996
rect 20656 11942 20658 11994
rect 20658 11942 20710 11994
rect 20710 11942 20712 11994
rect 20736 11942 20774 11994
rect 20774 11942 20786 11994
rect 20786 11942 20792 11994
rect 20816 11942 20838 11994
rect 20838 11942 20850 11994
rect 20850 11942 20872 11994
rect 20896 11942 20902 11994
rect 20902 11942 20914 11994
rect 20914 11942 20952 11994
rect 20976 11942 20978 11994
rect 20978 11942 21030 11994
rect 21030 11942 21032 11994
rect 20656 11940 20712 11942
rect 20736 11940 20792 11942
rect 20816 11940 20872 11942
rect 20896 11940 20952 11942
rect 20976 11940 21032 11942
rect 21086 11192 21142 11248
rect 20656 10906 20712 10908
rect 20736 10906 20792 10908
rect 20816 10906 20872 10908
rect 20896 10906 20952 10908
rect 20976 10906 21032 10908
rect 20656 10854 20658 10906
rect 20658 10854 20710 10906
rect 20710 10854 20712 10906
rect 20736 10854 20774 10906
rect 20774 10854 20786 10906
rect 20786 10854 20792 10906
rect 20816 10854 20838 10906
rect 20838 10854 20850 10906
rect 20850 10854 20872 10906
rect 20896 10854 20902 10906
rect 20902 10854 20914 10906
rect 20914 10854 20952 10906
rect 20976 10854 20978 10906
rect 20978 10854 21030 10906
rect 21030 10854 21032 10906
rect 20656 10852 20712 10854
rect 20736 10852 20792 10854
rect 20816 10852 20872 10854
rect 20896 10852 20952 10854
rect 20976 10852 21032 10854
rect 20656 9818 20712 9820
rect 20736 9818 20792 9820
rect 20816 9818 20872 9820
rect 20896 9818 20952 9820
rect 20976 9818 21032 9820
rect 20656 9766 20658 9818
rect 20658 9766 20710 9818
rect 20710 9766 20712 9818
rect 20736 9766 20774 9818
rect 20774 9766 20786 9818
rect 20786 9766 20792 9818
rect 20816 9766 20838 9818
rect 20838 9766 20850 9818
rect 20850 9766 20872 9818
rect 20896 9766 20902 9818
rect 20902 9766 20914 9818
rect 20914 9766 20952 9818
rect 20976 9766 20978 9818
rect 20978 9766 21030 9818
rect 21030 9766 21032 9818
rect 20656 9764 20712 9766
rect 20736 9764 20792 9766
rect 20816 9764 20872 9766
rect 20896 9764 20952 9766
rect 20976 9764 21032 9766
rect 21178 10240 21234 10296
rect 20810 9580 20866 9616
rect 20810 9560 20812 9580
rect 20812 9560 20864 9580
rect 20864 9560 20866 9580
rect 20074 9424 20130 9480
rect 19916 9274 19972 9276
rect 19996 9274 20052 9276
rect 20076 9274 20132 9276
rect 20156 9274 20212 9276
rect 20236 9274 20292 9276
rect 19916 9222 19918 9274
rect 19918 9222 19970 9274
rect 19970 9222 19972 9274
rect 19996 9222 20034 9274
rect 20034 9222 20046 9274
rect 20046 9222 20052 9274
rect 20076 9222 20098 9274
rect 20098 9222 20110 9274
rect 20110 9222 20132 9274
rect 20156 9222 20162 9274
rect 20162 9222 20174 9274
rect 20174 9222 20212 9274
rect 20236 9222 20238 9274
rect 20238 9222 20290 9274
rect 20290 9222 20292 9274
rect 19916 9220 19972 9222
rect 19996 9220 20052 9222
rect 20076 9220 20132 9222
rect 20156 9220 20212 9222
rect 20236 9220 20292 9222
rect 21270 10104 21326 10160
rect 21178 9560 21234 9616
rect 20656 8730 20712 8732
rect 20736 8730 20792 8732
rect 20816 8730 20872 8732
rect 20896 8730 20952 8732
rect 20976 8730 21032 8732
rect 20656 8678 20658 8730
rect 20658 8678 20710 8730
rect 20710 8678 20712 8730
rect 20736 8678 20774 8730
rect 20774 8678 20786 8730
rect 20786 8678 20792 8730
rect 20816 8678 20838 8730
rect 20838 8678 20850 8730
rect 20850 8678 20872 8730
rect 20896 8678 20902 8730
rect 20902 8678 20914 8730
rect 20914 8678 20952 8730
rect 20976 8678 20978 8730
rect 20978 8678 21030 8730
rect 21030 8678 21032 8730
rect 20656 8676 20712 8678
rect 20736 8676 20792 8678
rect 20816 8676 20872 8678
rect 20896 8676 20952 8678
rect 20976 8676 21032 8678
rect 19916 8186 19972 8188
rect 19996 8186 20052 8188
rect 20076 8186 20132 8188
rect 20156 8186 20212 8188
rect 20236 8186 20292 8188
rect 19916 8134 19918 8186
rect 19918 8134 19970 8186
rect 19970 8134 19972 8186
rect 19996 8134 20034 8186
rect 20034 8134 20046 8186
rect 20046 8134 20052 8186
rect 20076 8134 20098 8186
rect 20098 8134 20110 8186
rect 20110 8134 20132 8186
rect 20156 8134 20162 8186
rect 20162 8134 20174 8186
rect 20174 8134 20212 8186
rect 20236 8134 20238 8186
rect 20238 8134 20290 8186
rect 20290 8134 20292 8186
rect 19916 8132 19972 8134
rect 19996 8132 20052 8134
rect 20076 8132 20132 8134
rect 20156 8132 20212 8134
rect 20236 8132 20292 8134
rect 19916 7098 19972 7100
rect 19996 7098 20052 7100
rect 20076 7098 20132 7100
rect 20156 7098 20212 7100
rect 20236 7098 20292 7100
rect 19916 7046 19918 7098
rect 19918 7046 19970 7098
rect 19970 7046 19972 7098
rect 19996 7046 20034 7098
rect 20034 7046 20046 7098
rect 20046 7046 20052 7098
rect 20076 7046 20098 7098
rect 20098 7046 20110 7098
rect 20110 7046 20132 7098
rect 20156 7046 20162 7098
rect 20162 7046 20174 7098
rect 20174 7046 20212 7098
rect 20236 7046 20238 7098
rect 20238 7046 20290 7098
rect 20290 7046 20292 7098
rect 19916 7044 19972 7046
rect 19996 7044 20052 7046
rect 20076 7044 20132 7046
rect 20156 7044 20212 7046
rect 20236 7044 20292 7046
rect 19916 6010 19972 6012
rect 19996 6010 20052 6012
rect 20076 6010 20132 6012
rect 20156 6010 20212 6012
rect 20236 6010 20292 6012
rect 19916 5958 19918 6010
rect 19918 5958 19970 6010
rect 19970 5958 19972 6010
rect 19996 5958 20034 6010
rect 20034 5958 20046 6010
rect 20046 5958 20052 6010
rect 20076 5958 20098 6010
rect 20098 5958 20110 6010
rect 20110 5958 20132 6010
rect 20156 5958 20162 6010
rect 20162 5958 20174 6010
rect 20174 5958 20212 6010
rect 20236 5958 20238 6010
rect 20238 5958 20290 6010
rect 20290 5958 20292 6010
rect 19916 5956 19972 5958
rect 19996 5956 20052 5958
rect 20076 5956 20132 5958
rect 20156 5956 20212 5958
rect 20236 5956 20292 5958
rect 20656 7642 20712 7644
rect 20736 7642 20792 7644
rect 20816 7642 20872 7644
rect 20896 7642 20952 7644
rect 20976 7642 21032 7644
rect 20656 7590 20658 7642
rect 20658 7590 20710 7642
rect 20710 7590 20712 7642
rect 20736 7590 20774 7642
rect 20774 7590 20786 7642
rect 20786 7590 20792 7642
rect 20816 7590 20838 7642
rect 20838 7590 20850 7642
rect 20850 7590 20872 7642
rect 20896 7590 20902 7642
rect 20902 7590 20914 7642
rect 20914 7590 20952 7642
rect 20976 7590 20978 7642
rect 20978 7590 21030 7642
rect 21030 7590 21032 7642
rect 20656 7588 20712 7590
rect 20736 7588 20792 7590
rect 20816 7588 20872 7590
rect 20896 7588 20952 7590
rect 20976 7588 21032 7590
rect 21454 10240 21510 10296
rect 21362 9460 21364 9480
rect 21364 9460 21416 9480
rect 21416 9460 21418 9480
rect 21362 9424 21418 9460
rect 20656 6554 20712 6556
rect 20736 6554 20792 6556
rect 20816 6554 20872 6556
rect 20896 6554 20952 6556
rect 20976 6554 21032 6556
rect 20656 6502 20658 6554
rect 20658 6502 20710 6554
rect 20710 6502 20712 6554
rect 20736 6502 20774 6554
rect 20774 6502 20786 6554
rect 20786 6502 20792 6554
rect 20816 6502 20838 6554
rect 20838 6502 20850 6554
rect 20850 6502 20872 6554
rect 20896 6502 20902 6554
rect 20902 6502 20914 6554
rect 20914 6502 20952 6554
rect 20976 6502 20978 6554
rect 20978 6502 21030 6554
rect 21030 6502 21032 6554
rect 20656 6500 20712 6502
rect 20736 6500 20792 6502
rect 20816 6500 20872 6502
rect 20896 6500 20952 6502
rect 20976 6500 21032 6502
rect 21730 9560 21786 9616
rect 21638 9424 21694 9480
rect 20656 5466 20712 5468
rect 20736 5466 20792 5468
rect 20816 5466 20872 5468
rect 20896 5466 20952 5468
rect 20976 5466 21032 5468
rect 20656 5414 20658 5466
rect 20658 5414 20710 5466
rect 20710 5414 20712 5466
rect 20736 5414 20774 5466
rect 20774 5414 20786 5466
rect 20786 5414 20792 5466
rect 20816 5414 20838 5466
rect 20838 5414 20850 5466
rect 20850 5414 20872 5466
rect 20896 5414 20902 5466
rect 20902 5414 20914 5466
rect 20914 5414 20952 5466
rect 20976 5414 20978 5466
rect 20978 5414 21030 5466
rect 21030 5414 21032 5466
rect 20656 5412 20712 5414
rect 20736 5412 20792 5414
rect 20816 5412 20872 5414
rect 20896 5412 20952 5414
rect 20976 5412 21032 5414
rect 19916 4922 19972 4924
rect 19996 4922 20052 4924
rect 20076 4922 20132 4924
rect 20156 4922 20212 4924
rect 20236 4922 20292 4924
rect 19916 4870 19918 4922
rect 19918 4870 19970 4922
rect 19970 4870 19972 4922
rect 19996 4870 20034 4922
rect 20034 4870 20046 4922
rect 20046 4870 20052 4922
rect 20076 4870 20098 4922
rect 20098 4870 20110 4922
rect 20110 4870 20132 4922
rect 20156 4870 20162 4922
rect 20162 4870 20174 4922
rect 20174 4870 20212 4922
rect 20236 4870 20238 4922
rect 20238 4870 20290 4922
rect 20290 4870 20292 4922
rect 19916 4868 19972 4870
rect 19996 4868 20052 4870
rect 20076 4868 20132 4870
rect 20156 4868 20212 4870
rect 20236 4868 20292 4870
rect 22650 12280 22706 12336
rect 22466 10920 22522 10976
rect 22282 10104 22338 10160
rect 23294 16360 23350 16416
rect 23294 15680 23350 15736
rect 23386 14340 23442 14376
rect 23386 14320 23388 14340
rect 23388 14320 23440 14340
rect 23440 14320 23442 14340
rect 23386 13640 23442 13696
rect 23386 12960 23442 13016
rect 23202 11600 23258 11656
rect 23110 11192 23166 11248
rect 22742 10512 22798 10568
rect 23294 9444 23350 9480
rect 23294 9424 23296 9444
rect 23296 9424 23348 9444
rect 23348 9424 23350 9444
rect 20656 4378 20712 4380
rect 20736 4378 20792 4380
rect 20816 4378 20872 4380
rect 20896 4378 20952 4380
rect 20976 4378 21032 4380
rect 20656 4326 20658 4378
rect 20658 4326 20710 4378
rect 20710 4326 20712 4378
rect 20736 4326 20774 4378
rect 20774 4326 20786 4378
rect 20786 4326 20792 4378
rect 20816 4326 20838 4378
rect 20838 4326 20850 4378
rect 20850 4326 20872 4378
rect 20896 4326 20902 4378
rect 20902 4326 20914 4378
rect 20914 4326 20952 4378
rect 20976 4326 20978 4378
rect 20978 4326 21030 4378
rect 21030 4326 21032 4378
rect 20656 4324 20712 4326
rect 20736 4324 20792 4326
rect 20816 4324 20872 4326
rect 20896 4324 20952 4326
rect 20976 4324 21032 4326
rect 23018 8880 23074 8936
rect 23294 8200 23350 8256
rect 19916 3834 19972 3836
rect 19996 3834 20052 3836
rect 20076 3834 20132 3836
rect 20156 3834 20212 3836
rect 20236 3834 20292 3836
rect 19916 3782 19918 3834
rect 19918 3782 19970 3834
rect 19970 3782 19972 3834
rect 19996 3782 20034 3834
rect 20034 3782 20046 3834
rect 20046 3782 20052 3834
rect 20076 3782 20098 3834
rect 20098 3782 20110 3834
rect 20110 3782 20132 3834
rect 20156 3782 20162 3834
rect 20162 3782 20174 3834
rect 20174 3782 20212 3834
rect 20236 3782 20238 3834
rect 20238 3782 20290 3834
rect 20290 3782 20292 3834
rect 19916 3780 19972 3782
rect 19996 3780 20052 3782
rect 20076 3780 20132 3782
rect 20156 3780 20212 3782
rect 20236 3780 20292 3782
rect 20656 3290 20712 3292
rect 20736 3290 20792 3292
rect 20816 3290 20872 3292
rect 20896 3290 20952 3292
rect 20976 3290 21032 3292
rect 20656 3238 20658 3290
rect 20658 3238 20710 3290
rect 20710 3238 20712 3290
rect 20736 3238 20774 3290
rect 20774 3238 20786 3290
rect 20786 3238 20792 3290
rect 20816 3238 20838 3290
rect 20838 3238 20850 3290
rect 20850 3238 20872 3290
rect 20896 3238 20902 3290
rect 20902 3238 20914 3290
rect 20914 3238 20952 3290
rect 20976 3238 20978 3290
rect 20978 3238 21030 3290
rect 21030 3238 21032 3290
rect 20656 3236 20712 3238
rect 20736 3236 20792 3238
rect 20816 3236 20872 3238
rect 20896 3236 20952 3238
rect 20976 3236 21032 3238
rect 19916 2746 19972 2748
rect 19996 2746 20052 2748
rect 20076 2746 20132 2748
rect 20156 2746 20212 2748
rect 20236 2746 20292 2748
rect 19916 2694 19918 2746
rect 19918 2694 19970 2746
rect 19970 2694 19972 2746
rect 19996 2694 20034 2746
rect 20034 2694 20046 2746
rect 20046 2694 20052 2746
rect 20076 2694 20098 2746
rect 20098 2694 20110 2746
rect 20110 2694 20132 2746
rect 20156 2694 20162 2746
rect 20162 2694 20174 2746
rect 20174 2694 20212 2746
rect 20236 2694 20238 2746
rect 20238 2694 20290 2746
rect 20290 2694 20292 2746
rect 19916 2692 19972 2694
rect 19996 2692 20052 2694
rect 20076 2692 20132 2694
rect 20156 2692 20212 2694
rect 20236 2692 20292 2694
rect 14656 2202 14712 2204
rect 14736 2202 14792 2204
rect 14816 2202 14872 2204
rect 14896 2202 14952 2204
rect 14976 2202 15032 2204
rect 14656 2150 14658 2202
rect 14658 2150 14710 2202
rect 14710 2150 14712 2202
rect 14736 2150 14774 2202
rect 14774 2150 14786 2202
rect 14786 2150 14792 2202
rect 14816 2150 14838 2202
rect 14838 2150 14850 2202
rect 14850 2150 14872 2202
rect 14896 2150 14902 2202
rect 14902 2150 14914 2202
rect 14914 2150 14952 2202
rect 14976 2150 14978 2202
rect 14978 2150 15030 2202
rect 15030 2150 15032 2202
rect 14656 2148 14712 2150
rect 14736 2148 14792 2150
rect 14816 2148 14872 2150
rect 14896 2148 14952 2150
rect 14976 2148 15032 2150
rect 20656 2202 20712 2204
rect 20736 2202 20792 2204
rect 20816 2202 20872 2204
rect 20896 2202 20952 2204
rect 20976 2202 21032 2204
rect 20656 2150 20658 2202
rect 20658 2150 20710 2202
rect 20710 2150 20712 2202
rect 20736 2150 20774 2202
rect 20774 2150 20786 2202
rect 20786 2150 20792 2202
rect 20816 2150 20838 2202
rect 20838 2150 20850 2202
rect 20850 2150 20872 2202
rect 20896 2150 20902 2202
rect 20902 2150 20914 2202
rect 20914 2150 20952 2202
rect 20976 2150 20978 2202
rect 20978 2150 21030 2202
rect 21030 2150 21032 2202
rect 20656 2148 20712 2150
rect 20736 2148 20792 2150
rect 20816 2148 20872 2150
rect 20896 2148 20952 2150
rect 20976 2148 21032 2150
<< metal3 >>
rect 1906 24512 2302 24513
rect 1906 24448 1912 24512
rect 1976 24448 1992 24512
rect 2056 24448 2072 24512
rect 2136 24448 2152 24512
rect 2216 24448 2232 24512
rect 2296 24448 2302 24512
rect 1906 24447 2302 24448
rect 7906 24512 8302 24513
rect 7906 24448 7912 24512
rect 7976 24448 7992 24512
rect 8056 24448 8072 24512
rect 8136 24448 8152 24512
rect 8216 24448 8232 24512
rect 8296 24448 8302 24512
rect 7906 24447 8302 24448
rect 13906 24512 14302 24513
rect 13906 24448 13912 24512
rect 13976 24448 13992 24512
rect 14056 24448 14072 24512
rect 14136 24448 14152 24512
rect 14216 24448 14232 24512
rect 14296 24448 14302 24512
rect 13906 24447 14302 24448
rect 19906 24512 20302 24513
rect 19906 24448 19912 24512
rect 19976 24448 19992 24512
rect 20056 24448 20072 24512
rect 20136 24448 20152 24512
rect 20216 24448 20232 24512
rect 20296 24448 20302 24512
rect 19906 24447 20302 24448
rect 2646 23968 3042 23969
rect 2646 23904 2652 23968
rect 2716 23904 2732 23968
rect 2796 23904 2812 23968
rect 2876 23904 2892 23968
rect 2956 23904 2972 23968
rect 3036 23904 3042 23968
rect 2646 23903 3042 23904
rect 8646 23968 9042 23969
rect 8646 23904 8652 23968
rect 8716 23904 8732 23968
rect 8796 23904 8812 23968
rect 8876 23904 8892 23968
rect 8956 23904 8972 23968
rect 9036 23904 9042 23968
rect 8646 23903 9042 23904
rect 14646 23968 15042 23969
rect 14646 23904 14652 23968
rect 14716 23904 14732 23968
rect 14796 23904 14812 23968
rect 14876 23904 14892 23968
rect 14956 23904 14972 23968
rect 15036 23904 15042 23968
rect 14646 23903 15042 23904
rect 20646 23968 21042 23969
rect 20646 23904 20652 23968
rect 20716 23904 20732 23968
rect 20796 23904 20812 23968
rect 20876 23904 20892 23968
rect 20956 23904 20972 23968
rect 21036 23904 21042 23968
rect 20646 23903 21042 23904
rect 1906 23424 2302 23425
rect 1906 23360 1912 23424
rect 1976 23360 1992 23424
rect 2056 23360 2072 23424
rect 2136 23360 2152 23424
rect 2216 23360 2232 23424
rect 2296 23360 2302 23424
rect 1906 23359 2302 23360
rect 7906 23424 8302 23425
rect 7906 23360 7912 23424
rect 7976 23360 7992 23424
rect 8056 23360 8072 23424
rect 8136 23360 8152 23424
rect 8216 23360 8232 23424
rect 8296 23360 8302 23424
rect 7906 23359 8302 23360
rect 13906 23424 14302 23425
rect 13906 23360 13912 23424
rect 13976 23360 13992 23424
rect 14056 23360 14072 23424
rect 14136 23360 14152 23424
rect 14216 23360 14232 23424
rect 14296 23360 14302 23424
rect 13906 23359 14302 23360
rect 19906 23424 20302 23425
rect 19906 23360 19912 23424
rect 19976 23360 19992 23424
rect 20056 23360 20072 23424
rect 20136 23360 20152 23424
rect 20216 23360 20232 23424
rect 20296 23360 20302 23424
rect 19906 23359 20302 23360
rect 2646 22880 3042 22881
rect 2646 22816 2652 22880
rect 2716 22816 2732 22880
rect 2796 22816 2812 22880
rect 2876 22816 2892 22880
rect 2956 22816 2972 22880
rect 3036 22816 3042 22880
rect 2646 22815 3042 22816
rect 8646 22880 9042 22881
rect 8646 22816 8652 22880
rect 8716 22816 8732 22880
rect 8796 22816 8812 22880
rect 8876 22816 8892 22880
rect 8956 22816 8972 22880
rect 9036 22816 9042 22880
rect 8646 22815 9042 22816
rect 14646 22880 15042 22881
rect 14646 22816 14652 22880
rect 14716 22816 14732 22880
rect 14796 22816 14812 22880
rect 14876 22816 14892 22880
rect 14956 22816 14972 22880
rect 15036 22816 15042 22880
rect 14646 22815 15042 22816
rect 20646 22880 21042 22881
rect 20646 22816 20652 22880
rect 20716 22816 20732 22880
rect 20796 22816 20812 22880
rect 20876 22816 20892 22880
rect 20956 22816 20972 22880
rect 21036 22816 21042 22880
rect 20646 22815 21042 22816
rect 1906 22336 2302 22337
rect 1906 22272 1912 22336
rect 1976 22272 1992 22336
rect 2056 22272 2072 22336
rect 2136 22272 2152 22336
rect 2216 22272 2232 22336
rect 2296 22272 2302 22336
rect 1906 22271 2302 22272
rect 7906 22336 8302 22337
rect 7906 22272 7912 22336
rect 7976 22272 7992 22336
rect 8056 22272 8072 22336
rect 8136 22272 8152 22336
rect 8216 22272 8232 22336
rect 8296 22272 8302 22336
rect 7906 22271 8302 22272
rect 13906 22336 14302 22337
rect 13906 22272 13912 22336
rect 13976 22272 13992 22336
rect 14056 22272 14072 22336
rect 14136 22272 14152 22336
rect 14216 22272 14232 22336
rect 14296 22272 14302 22336
rect 13906 22271 14302 22272
rect 19906 22336 20302 22337
rect 19906 22272 19912 22336
rect 19976 22272 19992 22336
rect 20056 22272 20072 22336
rect 20136 22272 20152 22336
rect 20216 22272 20232 22336
rect 20296 22272 20302 22336
rect 19906 22271 20302 22272
rect 2646 21792 3042 21793
rect 2646 21728 2652 21792
rect 2716 21728 2732 21792
rect 2796 21728 2812 21792
rect 2876 21728 2892 21792
rect 2956 21728 2972 21792
rect 3036 21728 3042 21792
rect 2646 21727 3042 21728
rect 8646 21792 9042 21793
rect 8646 21728 8652 21792
rect 8716 21728 8732 21792
rect 8796 21728 8812 21792
rect 8876 21728 8892 21792
rect 8956 21728 8972 21792
rect 9036 21728 9042 21792
rect 8646 21727 9042 21728
rect 14646 21792 15042 21793
rect 14646 21728 14652 21792
rect 14716 21728 14732 21792
rect 14796 21728 14812 21792
rect 14876 21728 14892 21792
rect 14956 21728 14972 21792
rect 15036 21728 15042 21792
rect 14646 21727 15042 21728
rect 20646 21792 21042 21793
rect 20646 21728 20652 21792
rect 20716 21728 20732 21792
rect 20796 21728 20812 21792
rect 20876 21728 20892 21792
rect 20956 21728 20972 21792
rect 21036 21728 21042 21792
rect 20646 21727 21042 21728
rect 1906 21248 2302 21249
rect 1906 21184 1912 21248
rect 1976 21184 1992 21248
rect 2056 21184 2072 21248
rect 2136 21184 2152 21248
rect 2216 21184 2232 21248
rect 2296 21184 2302 21248
rect 1906 21183 2302 21184
rect 7906 21248 8302 21249
rect 7906 21184 7912 21248
rect 7976 21184 7992 21248
rect 8056 21184 8072 21248
rect 8136 21184 8152 21248
rect 8216 21184 8232 21248
rect 8296 21184 8302 21248
rect 7906 21183 8302 21184
rect 13906 21248 14302 21249
rect 13906 21184 13912 21248
rect 13976 21184 13992 21248
rect 14056 21184 14072 21248
rect 14136 21184 14152 21248
rect 14216 21184 14232 21248
rect 14296 21184 14302 21248
rect 13906 21183 14302 21184
rect 19906 21248 20302 21249
rect 19906 21184 19912 21248
rect 19976 21184 19992 21248
rect 20056 21184 20072 21248
rect 20136 21184 20152 21248
rect 20216 21184 20232 21248
rect 20296 21184 20302 21248
rect 19906 21183 20302 21184
rect 2646 20704 3042 20705
rect 2646 20640 2652 20704
rect 2716 20640 2732 20704
rect 2796 20640 2812 20704
rect 2876 20640 2892 20704
rect 2956 20640 2972 20704
rect 3036 20640 3042 20704
rect 2646 20639 3042 20640
rect 8646 20704 9042 20705
rect 8646 20640 8652 20704
rect 8716 20640 8732 20704
rect 8796 20640 8812 20704
rect 8876 20640 8892 20704
rect 8956 20640 8972 20704
rect 9036 20640 9042 20704
rect 8646 20639 9042 20640
rect 14646 20704 15042 20705
rect 14646 20640 14652 20704
rect 14716 20640 14732 20704
rect 14796 20640 14812 20704
rect 14876 20640 14892 20704
rect 14956 20640 14972 20704
rect 15036 20640 15042 20704
rect 14646 20639 15042 20640
rect 20646 20704 21042 20705
rect 20646 20640 20652 20704
rect 20716 20640 20732 20704
rect 20796 20640 20812 20704
rect 20876 20640 20892 20704
rect 20956 20640 20972 20704
rect 21036 20640 21042 20704
rect 20646 20639 21042 20640
rect 1906 20160 2302 20161
rect 1906 20096 1912 20160
rect 1976 20096 1992 20160
rect 2056 20096 2072 20160
rect 2136 20096 2152 20160
rect 2216 20096 2232 20160
rect 2296 20096 2302 20160
rect 1906 20095 2302 20096
rect 7906 20160 8302 20161
rect 7906 20096 7912 20160
rect 7976 20096 7992 20160
rect 8056 20096 8072 20160
rect 8136 20096 8152 20160
rect 8216 20096 8232 20160
rect 8296 20096 8302 20160
rect 7906 20095 8302 20096
rect 13906 20160 14302 20161
rect 13906 20096 13912 20160
rect 13976 20096 13992 20160
rect 14056 20096 14072 20160
rect 14136 20096 14152 20160
rect 14216 20096 14232 20160
rect 14296 20096 14302 20160
rect 13906 20095 14302 20096
rect 19906 20160 20302 20161
rect 19906 20096 19912 20160
rect 19976 20096 19992 20160
rect 20056 20096 20072 20160
rect 20136 20096 20152 20160
rect 20216 20096 20232 20160
rect 20296 20096 20302 20160
rect 19906 20095 20302 20096
rect 0 19818 800 19848
rect 3785 19818 3851 19821
rect 0 19816 3851 19818
rect 0 19760 3790 19816
rect 3846 19760 3851 19816
rect 0 19758 3851 19760
rect 0 19728 800 19758
rect 3785 19755 3851 19758
rect 2646 19616 3042 19617
rect 2646 19552 2652 19616
rect 2716 19552 2732 19616
rect 2796 19552 2812 19616
rect 2876 19552 2892 19616
rect 2956 19552 2972 19616
rect 3036 19552 3042 19616
rect 2646 19551 3042 19552
rect 8646 19616 9042 19617
rect 8646 19552 8652 19616
rect 8716 19552 8732 19616
rect 8796 19552 8812 19616
rect 8876 19552 8892 19616
rect 8956 19552 8972 19616
rect 9036 19552 9042 19616
rect 8646 19551 9042 19552
rect 14646 19616 15042 19617
rect 14646 19552 14652 19616
rect 14716 19552 14732 19616
rect 14796 19552 14812 19616
rect 14876 19552 14892 19616
rect 14956 19552 14972 19616
rect 15036 19552 15042 19616
rect 14646 19551 15042 19552
rect 20646 19616 21042 19617
rect 20646 19552 20652 19616
rect 20716 19552 20732 19616
rect 20796 19552 20812 19616
rect 20876 19552 20892 19616
rect 20956 19552 20972 19616
rect 21036 19552 21042 19616
rect 20646 19551 21042 19552
rect 14917 19410 14983 19413
rect 15561 19410 15627 19413
rect 14917 19408 15627 19410
rect 14917 19352 14922 19408
rect 14978 19352 15566 19408
rect 15622 19352 15627 19408
rect 14917 19350 15627 19352
rect 14917 19347 14983 19350
rect 15561 19347 15627 19350
rect 23289 19138 23355 19141
rect 24200 19138 25000 19168
rect 23289 19136 25000 19138
rect 23289 19080 23294 19136
rect 23350 19080 25000 19136
rect 23289 19078 25000 19080
rect 23289 19075 23355 19078
rect 1906 19072 2302 19073
rect 1906 19008 1912 19072
rect 1976 19008 1992 19072
rect 2056 19008 2072 19072
rect 2136 19008 2152 19072
rect 2216 19008 2232 19072
rect 2296 19008 2302 19072
rect 1906 19007 2302 19008
rect 7906 19072 8302 19073
rect 7906 19008 7912 19072
rect 7976 19008 7992 19072
rect 8056 19008 8072 19072
rect 8136 19008 8152 19072
rect 8216 19008 8232 19072
rect 8296 19008 8302 19072
rect 7906 19007 8302 19008
rect 13906 19072 14302 19073
rect 13906 19008 13912 19072
rect 13976 19008 13992 19072
rect 14056 19008 14072 19072
rect 14136 19008 14152 19072
rect 14216 19008 14232 19072
rect 14296 19008 14302 19072
rect 13906 19007 14302 19008
rect 19906 19072 20302 19073
rect 19906 19008 19912 19072
rect 19976 19008 19992 19072
rect 20056 19008 20072 19072
rect 20136 19008 20152 19072
rect 20216 19008 20232 19072
rect 20296 19008 20302 19072
rect 24200 19048 25000 19078
rect 19906 19007 20302 19008
rect 2646 18528 3042 18529
rect 2646 18464 2652 18528
rect 2716 18464 2732 18528
rect 2796 18464 2812 18528
rect 2876 18464 2892 18528
rect 2956 18464 2972 18528
rect 3036 18464 3042 18528
rect 2646 18463 3042 18464
rect 8646 18528 9042 18529
rect 8646 18464 8652 18528
rect 8716 18464 8732 18528
rect 8796 18464 8812 18528
rect 8876 18464 8892 18528
rect 8956 18464 8972 18528
rect 9036 18464 9042 18528
rect 8646 18463 9042 18464
rect 14646 18528 15042 18529
rect 14646 18464 14652 18528
rect 14716 18464 14732 18528
rect 14796 18464 14812 18528
rect 14876 18464 14892 18528
rect 14956 18464 14972 18528
rect 15036 18464 15042 18528
rect 14646 18463 15042 18464
rect 20646 18528 21042 18529
rect 20646 18464 20652 18528
rect 20716 18464 20732 18528
rect 20796 18464 20812 18528
rect 20876 18464 20892 18528
rect 20956 18464 20972 18528
rect 21036 18464 21042 18528
rect 20646 18463 21042 18464
rect 23289 18458 23355 18461
rect 24200 18458 25000 18488
rect 23289 18456 25000 18458
rect 23289 18400 23294 18456
rect 23350 18400 25000 18456
rect 23289 18398 25000 18400
rect 23289 18395 23355 18398
rect 24200 18368 25000 18398
rect 1906 17984 2302 17985
rect 1906 17920 1912 17984
rect 1976 17920 1992 17984
rect 2056 17920 2072 17984
rect 2136 17920 2152 17984
rect 2216 17920 2232 17984
rect 2296 17920 2302 17984
rect 1906 17919 2302 17920
rect 7906 17984 8302 17985
rect 7906 17920 7912 17984
rect 7976 17920 7992 17984
rect 8056 17920 8072 17984
rect 8136 17920 8152 17984
rect 8216 17920 8232 17984
rect 8296 17920 8302 17984
rect 7906 17919 8302 17920
rect 13906 17984 14302 17985
rect 13906 17920 13912 17984
rect 13976 17920 13992 17984
rect 14056 17920 14072 17984
rect 14136 17920 14152 17984
rect 14216 17920 14232 17984
rect 14296 17920 14302 17984
rect 13906 17919 14302 17920
rect 19906 17984 20302 17985
rect 19906 17920 19912 17984
rect 19976 17920 19992 17984
rect 20056 17920 20072 17984
rect 20136 17920 20152 17984
rect 20216 17920 20232 17984
rect 20296 17920 20302 17984
rect 19906 17919 20302 17920
rect 5349 17778 5415 17781
rect 10133 17778 10199 17781
rect 5349 17776 10199 17778
rect 5349 17720 5354 17776
rect 5410 17720 10138 17776
rect 10194 17720 10199 17776
rect 5349 17718 10199 17720
rect 5349 17715 5415 17718
rect 10133 17715 10199 17718
rect 2646 17440 3042 17441
rect 2646 17376 2652 17440
rect 2716 17376 2732 17440
rect 2796 17376 2812 17440
rect 2876 17376 2892 17440
rect 2956 17376 2972 17440
rect 3036 17376 3042 17440
rect 2646 17375 3042 17376
rect 8646 17440 9042 17441
rect 8646 17376 8652 17440
rect 8716 17376 8732 17440
rect 8796 17376 8812 17440
rect 8876 17376 8892 17440
rect 8956 17376 8972 17440
rect 9036 17376 9042 17440
rect 8646 17375 9042 17376
rect 14646 17440 15042 17441
rect 14646 17376 14652 17440
rect 14716 17376 14732 17440
rect 14796 17376 14812 17440
rect 14876 17376 14892 17440
rect 14956 17376 14972 17440
rect 15036 17376 15042 17440
rect 14646 17375 15042 17376
rect 20646 17440 21042 17441
rect 20646 17376 20652 17440
rect 20716 17376 20732 17440
rect 20796 17376 20812 17440
rect 20876 17376 20892 17440
rect 20956 17376 20972 17440
rect 21036 17376 21042 17440
rect 20646 17375 21042 17376
rect 0 17098 800 17128
rect 933 17098 999 17101
rect 0 17096 999 17098
rect 0 17040 938 17096
rect 994 17040 999 17096
rect 0 17038 999 17040
rect 0 17008 800 17038
rect 933 17035 999 17038
rect 3417 17098 3483 17101
rect 8661 17098 8727 17101
rect 3417 17096 8727 17098
rect 3417 17040 3422 17096
rect 3478 17040 8666 17096
rect 8722 17040 8727 17096
rect 3417 17038 8727 17040
rect 3417 17035 3483 17038
rect 8661 17035 8727 17038
rect 1906 16896 2302 16897
rect 1906 16832 1912 16896
rect 1976 16832 1992 16896
rect 2056 16832 2072 16896
rect 2136 16832 2152 16896
rect 2216 16832 2232 16896
rect 2296 16832 2302 16896
rect 1906 16831 2302 16832
rect 7906 16896 8302 16897
rect 7906 16832 7912 16896
rect 7976 16832 7992 16896
rect 8056 16832 8072 16896
rect 8136 16832 8152 16896
rect 8216 16832 8232 16896
rect 8296 16832 8302 16896
rect 7906 16831 8302 16832
rect 13906 16896 14302 16897
rect 13906 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14152 16896
rect 14216 16832 14232 16896
rect 14296 16832 14302 16896
rect 13906 16831 14302 16832
rect 19906 16896 20302 16897
rect 19906 16832 19912 16896
rect 19976 16832 19992 16896
rect 20056 16832 20072 16896
rect 20136 16832 20152 16896
rect 20216 16832 20232 16896
rect 20296 16832 20302 16896
rect 19906 16831 20302 16832
rect 3877 16690 3943 16693
rect 9029 16690 9095 16693
rect 3877 16688 9095 16690
rect 3877 16632 3882 16688
rect 3938 16632 9034 16688
rect 9090 16632 9095 16688
rect 3877 16630 9095 16632
rect 3877 16627 3943 16630
rect 9029 16627 9095 16630
rect 23289 16418 23355 16421
rect 24200 16418 25000 16448
rect 23289 16416 25000 16418
rect 23289 16360 23294 16416
rect 23350 16360 25000 16416
rect 23289 16358 25000 16360
rect 23289 16355 23355 16358
rect 2646 16352 3042 16353
rect 2646 16288 2652 16352
rect 2716 16288 2732 16352
rect 2796 16288 2812 16352
rect 2876 16288 2892 16352
rect 2956 16288 2972 16352
rect 3036 16288 3042 16352
rect 2646 16287 3042 16288
rect 8646 16352 9042 16353
rect 8646 16288 8652 16352
rect 8716 16288 8732 16352
rect 8796 16288 8812 16352
rect 8876 16288 8892 16352
rect 8956 16288 8972 16352
rect 9036 16288 9042 16352
rect 8646 16287 9042 16288
rect 14646 16352 15042 16353
rect 14646 16288 14652 16352
rect 14716 16288 14732 16352
rect 14796 16288 14812 16352
rect 14876 16288 14892 16352
rect 14956 16288 14972 16352
rect 15036 16288 15042 16352
rect 14646 16287 15042 16288
rect 20646 16352 21042 16353
rect 20646 16288 20652 16352
rect 20716 16288 20732 16352
rect 20796 16288 20812 16352
rect 20876 16288 20892 16352
rect 20956 16288 20972 16352
rect 21036 16288 21042 16352
rect 24200 16328 25000 16358
rect 20646 16287 21042 16288
rect 3601 16146 3667 16149
rect 9121 16146 9187 16149
rect 3601 16144 9187 16146
rect 3601 16088 3606 16144
rect 3662 16088 9126 16144
rect 9182 16088 9187 16144
rect 3601 16086 9187 16088
rect 3601 16083 3667 16086
rect 9121 16083 9187 16086
rect 1853 16010 1919 16013
rect 5349 16010 5415 16013
rect 8293 16010 8359 16013
rect 1853 16008 5415 16010
rect 1853 15952 1858 16008
rect 1914 15952 5354 16008
rect 5410 15952 5415 16008
rect 1853 15950 5415 15952
rect 1853 15947 1919 15950
rect 5349 15947 5415 15950
rect 5582 16008 8359 16010
rect 5582 15952 8298 16008
rect 8354 15952 8359 16008
rect 5582 15950 8359 15952
rect 1906 15808 2302 15809
rect 0 15738 800 15768
rect 1906 15744 1912 15808
rect 1976 15744 1992 15808
rect 2056 15744 2072 15808
rect 2136 15744 2152 15808
rect 2216 15744 2232 15808
rect 2296 15744 2302 15808
rect 1906 15743 2302 15744
rect 933 15738 999 15741
rect 5582 15738 5642 15950
rect 8293 15947 8359 15950
rect 7906 15808 8302 15809
rect 7906 15744 7912 15808
rect 7976 15744 7992 15808
rect 8056 15744 8072 15808
rect 8136 15744 8152 15808
rect 8216 15744 8232 15808
rect 8296 15744 8302 15808
rect 7906 15743 8302 15744
rect 13906 15808 14302 15809
rect 13906 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14152 15808
rect 14216 15744 14232 15808
rect 14296 15744 14302 15808
rect 13906 15743 14302 15744
rect 19906 15808 20302 15809
rect 19906 15744 19912 15808
rect 19976 15744 19992 15808
rect 20056 15744 20072 15808
rect 20136 15744 20152 15808
rect 20216 15744 20232 15808
rect 20296 15744 20302 15808
rect 19906 15743 20302 15744
rect 0 15736 999 15738
rect 0 15680 938 15736
rect 994 15680 999 15736
rect 0 15678 999 15680
rect 0 15648 800 15678
rect 933 15675 999 15678
rect 2730 15678 5642 15738
rect 23289 15738 23355 15741
rect 24200 15738 25000 15768
rect 23289 15736 25000 15738
rect 23289 15680 23294 15736
rect 23350 15680 25000 15736
rect 23289 15678 25000 15680
rect 2221 15602 2287 15605
rect 2730 15602 2790 15678
rect 23289 15675 23355 15678
rect 24200 15648 25000 15678
rect 2221 15600 2790 15602
rect 2221 15544 2226 15600
rect 2282 15544 2790 15600
rect 2221 15542 2790 15544
rect 3601 15602 3667 15605
rect 4797 15602 4863 15605
rect 3601 15600 4863 15602
rect 3601 15544 3606 15600
rect 3662 15544 4802 15600
rect 4858 15544 4863 15600
rect 3601 15542 4863 15544
rect 2221 15539 2287 15542
rect 3601 15539 3667 15542
rect 4797 15539 4863 15542
rect 2589 15466 2655 15469
rect 4245 15466 4311 15469
rect 2589 15464 4311 15466
rect 2589 15408 2594 15464
rect 2650 15408 4250 15464
rect 4306 15408 4311 15464
rect 2589 15406 4311 15408
rect 2589 15403 2655 15406
rect 4245 15403 4311 15406
rect 2646 15264 3042 15265
rect 2646 15200 2652 15264
rect 2716 15200 2732 15264
rect 2796 15200 2812 15264
rect 2876 15200 2892 15264
rect 2956 15200 2972 15264
rect 3036 15200 3042 15264
rect 2646 15199 3042 15200
rect 8646 15264 9042 15265
rect 8646 15200 8652 15264
rect 8716 15200 8732 15264
rect 8796 15200 8812 15264
rect 8876 15200 8892 15264
rect 8956 15200 8972 15264
rect 9036 15200 9042 15264
rect 8646 15199 9042 15200
rect 14646 15264 15042 15265
rect 14646 15200 14652 15264
rect 14716 15200 14732 15264
rect 14796 15200 14812 15264
rect 14876 15200 14892 15264
rect 14956 15200 14972 15264
rect 15036 15200 15042 15264
rect 14646 15199 15042 15200
rect 20646 15264 21042 15265
rect 20646 15200 20652 15264
rect 20716 15200 20732 15264
rect 20796 15200 20812 15264
rect 20876 15200 20892 15264
rect 20956 15200 20972 15264
rect 21036 15200 21042 15264
rect 20646 15199 21042 15200
rect 1906 14720 2302 14721
rect 1906 14656 1912 14720
rect 1976 14656 1992 14720
rect 2056 14656 2072 14720
rect 2136 14656 2152 14720
rect 2216 14656 2232 14720
rect 2296 14656 2302 14720
rect 1906 14655 2302 14656
rect 7906 14720 8302 14721
rect 7906 14656 7912 14720
rect 7976 14656 7992 14720
rect 8056 14656 8072 14720
rect 8136 14656 8152 14720
rect 8216 14656 8232 14720
rect 8296 14656 8302 14720
rect 7906 14655 8302 14656
rect 13906 14720 14302 14721
rect 13906 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14152 14720
rect 14216 14656 14232 14720
rect 14296 14656 14302 14720
rect 13906 14655 14302 14656
rect 19906 14720 20302 14721
rect 19906 14656 19912 14720
rect 19976 14656 19992 14720
rect 20056 14656 20072 14720
rect 20136 14656 20152 14720
rect 20216 14656 20232 14720
rect 20296 14656 20302 14720
rect 19906 14655 20302 14656
rect 23381 14378 23447 14381
rect 24200 14378 25000 14408
rect 23381 14376 25000 14378
rect 23381 14320 23386 14376
rect 23442 14320 25000 14376
rect 23381 14318 25000 14320
rect 23381 14315 23447 14318
rect 24200 14288 25000 14318
rect 2646 14176 3042 14177
rect 2646 14112 2652 14176
rect 2716 14112 2732 14176
rect 2796 14112 2812 14176
rect 2876 14112 2892 14176
rect 2956 14112 2972 14176
rect 3036 14112 3042 14176
rect 2646 14111 3042 14112
rect 8646 14176 9042 14177
rect 8646 14112 8652 14176
rect 8716 14112 8732 14176
rect 8796 14112 8812 14176
rect 8876 14112 8892 14176
rect 8956 14112 8972 14176
rect 9036 14112 9042 14176
rect 8646 14111 9042 14112
rect 14646 14176 15042 14177
rect 14646 14112 14652 14176
rect 14716 14112 14732 14176
rect 14796 14112 14812 14176
rect 14876 14112 14892 14176
rect 14956 14112 14972 14176
rect 15036 14112 15042 14176
rect 14646 14111 15042 14112
rect 20646 14176 21042 14177
rect 20646 14112 20652 14176
rect 20716 14112 20732 14176
rect 20796 14112 20812 14176
rect 20876 14112 20892 14176
rect 20956 14112 20972 14176
rect 21036 14112 21042 14176
rect 20646 14111 21042 14112
rect 0 13698 800 13728
rect 933 13698 999 13701
rect 0 13696 999 13698
rect 0 13640 938 13696
rect 994 13640 999 13696
rect 0 13638 999 13640
rect 0 13608 800 13638
rect 933 13635 999 13638
rect 23381 13698 23447 13701
rect 24200 13698 25000 13728
rect 23381 13696 25000 13698
rect 23381 13640 23386 13696
rect 23442 13640 25000 13696
rect 23381 13638 25000 13640
rect 23381 13635 23447 13638
rect 1906 13632 2302 13633
rect 1906 13568 1912 13632
rect 1976 13568 1992 13632
rect 2056 13568 2072 13632
rect 2136 13568 2152 13632
rect 2216 13568 2232 13632
rect 2296 13568 2302 13632
rect 1906 13567 2302 13568
rect 7906 13632 8302 13633
rect 7906 13568 7912 13632
rect 7976 13568 7992 13632
rect 8056 13568 8072 13632
rect 8136 13568 8152 13632
rect 8216 13568 8232 13632
rect 8296 13568 8302 13632
rect 7906 13567 8302 13568
rect 13906 13632 14302 13633
rect 13906 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14152 13632
rect 14216 13568 14232 13632
rect 14296 13568 14302 13632
rect 13906 13567 14302 13568
rect 19906 13632 20302 13633
rect 19906 13568 19912 13632
rect 19976 13568 19992 13632
rect 20056 13568 20072 13632
rect 20136 13568 20152 13632
rect 20216 13568 20232 13632
rect 20296 13568 20302 13632
rect 24200 13608 25000 13638
rect 19906 13567 20302 13568
rect 3785 13426 3851 13429
rect 11605 13426 11671 13429
rect 3785 13424 11671 13426
rect 3785 13368 3790 13424
rect 3846 13368 11610 13424
rect 11666 13368 11671 13424
rect 3785 13366 11671 13368
rect 3785 13363 3851 13366
rect 11605 13363 11671 13366
rect 14365 13426 14431 13429
rect 21541 13426 21607 13429
rect 14365 13424 21607 13426
rect 14365 13368 14370 13424
rect 14426 13368 21546 13424
rect 21602 13368 21607 13424
rect 14365 13366 21607 13368
rect 14365 13363 14431 13366
rect 21541 13363 21607 13366
rect 1301 13154 1367 13157
rect 936 13152 1367 13154
rect 936 13096 1306 13152
rect 1362 13096 1367 13152
rect 936 13094 1367 13096
rect 0 13018 800 13048
rect 936 13018 996 13094
rect 1301 13091 1367 13094
rect 2646 13088 3042 13089
rect 2646 13024 2652 13088
rect 2716 13024 2732 13088
rect 2796 13024 2812 13088
rect 2876 13024 2892 13088
rect 2956 13024 2972 13088
rect 3036 13024 3042 13088
rect 2646 13023 3042 13024
rect 8646 13088 9042 13089
rect 8646 13024 8652 13088
rect 8716 13024 8732 13088
rect 8796 13024 8812 13088
rect 8876 13024 8892 13088
rect 8956 13024 8972 13088
rect 9036 13024 9042 13088
rect 8646 13023 9042 13024
rect 14646 13088 15042 13089
rect 14646 13024 14652 13088
rect 14716 13024 14732 13088
rect 14796 13024 14812 13088
rect 14876 13024 14892 13088
rect 14956 13024 14972 13088
rect 15036 13024 15042 13088
rect 14646 13023 15042 13024
rect 20646 13088 21042 13089
rect 20646 13024 20652 13088
rect 20716 13024 20732 13088
rect 20796 13024 20812 13088
rect 20876 13024 20892 13088
rect 20956 13024 20972 13088
rect 21036 13024 21042 13088
rect 20646 13023 21042 13024
rect 0 12958 996 13018
rect 23381 13018 23447 13021
rect 24200 13018 25000 13048
rect 23381 13016 25000 13018
rect 23381 12960 23386 13016
rect 23442 12960 25000 13016
rect 23381 12958 25000 12960
rect 0 12928 800 12958
rect 23381 12955 23447 12958
rect 24200 12928 25000 12958
rect 3785 12882 3851 12885
rect 8385 12882 8451 12885
rect 3785 12880 8451 12882
rect 3785 12824 3790 12880
rect 3846 12824 8390 12880
rect 8446 12824 8451 12880
rect 3785 12822 8451 12824
rect 3785 12819 3851 12822
rect 8385 12819 8451 12822
rect 9397 12748 9463 12749
rect 9397 12744 9444 12748
rect 9508 12746 9514 12748
rect 14273 12746 14339 12749
rect 17217 12746 17283 12749
rect 9397 12688 9402 12744
rect 9397 12684 9444 12688
rect 9508 12686 9554 12746
rect 14273 12744 17283 12746
rect 14273 12688 14278 12744
rect 14334 12688 17222 12744
rect 17278 12688 17283 12744
rect 14273 12686 17283 12688
rect 9508 12684 9514 12686
rect 9397 12683 9463 12684
rect 14273 12683 14339 12686
rect 17217 12683 17283 12686
rect 9397 12610 9463 12613
rect 9765 12610 9831 12613
rect 9397 12608 9831 12610
rect 9397 12552 9402 12608
rect 9458 12552 9770 12608
rect 9826 12552 9831 12608
rect 9397 12550 9831 12552
rect 9397 12547 9463 12550
rect 9765 12547 9831 12550
rect 1906 12544 2302 12545
rect 1906 12480 1912 12544
rect 1976 12480 1992 12544
rect 2056 12480 2072 12544
rect 2136 12480 2152 12544
rect 2216 12480 2232 12544
rect 2296 12480 2302 12544
rect 1906 12479 2302 12480
rect 7906 12544 8302 12545
rect 7906 12480 7912 12544
rect 7976 12480 7992 12544
rect 8056 12480 8072 12544
rect 8136 12480 8152 12544
rect 8216 12480 8232 12544
rect 8296 12480 8302 12544
rect 7906 12479 8302 12480
rect 13906 12544 14302 12545
rect 13906 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14152 12544
rect 14216 12480 14232 12544
rect 14296 12480 14302 12544
rect 13906 12479 14302 12480
rect 19906 12544 20302 12545
rect 19906 12480 19912 12544
rect 19976 12480 19992 12544
rect 20056 12480 20072 12544
rect 20136 12480 20152 12544
rect 20216 12480 20232 12544
rect 20296 12480 20302 12544
rect 19906 12479 20302 12480
rect 0 12338 800 12368
rect 933 12338 999 12341
rect 0 12336 999 12338
rect 0 12280 938 12336
rect 994 12280 999 12336
rect 0 12278 999 12280
rect 0 12248 800 12278
rect 933 12275 999 12278
rect 22645 12338 22711 12341
rect 24200 12338 25000 12368
rect 22645 12336 25000 12338
rect 22645 12280 22650 12336
rect 22706 12280 25000 12336
rect 22645 12278 25000 12280
rect 22645 12275 22711 12278
rect 24200 12248 25000 12278
rect 2646 12000 3042 12001
rect 2646 11936 2652 12000
rect 2716 11936 2732 12000
rect 2796 11936 2812 12000
rect 2876 11936 2892 12000
rect 2956 11936 2972 12000
rect 3036 11936 3042 12000
rect 2646 11935 3042 11936
rect 8646 12000 9042 12001
rect 8646 11936 8652 12000
rect 8716 11936 8732 12000
rect 8796 11936 8812 12000
rect 8876 11936 8892 12000
rect 8956 11936 8972 12000
rect 9036 11936 9042 12000
rect 8646 11935 9042 11936
rect 14646 12000 15042 12001
rect 14646 11936 14652 12000
rect 14716 11936 14732 12000
rect 14796 11936 14812 12000
rect 14876 11936 14892 12000
rect 14956 11936 14972 12000
rect 15036 11936 15042 12000
rect 14646 11935 15042 11936
rect 20646 12000 21042 12001
rect 20646 11936 20652 12000
rect 20716 11936 20732 12000
rect 20796 11936 20812 12000
rect 20876 11936 20892 12000
rect 20956 11936 20972 12000
rect 21036 11936 21042 12000
rect 20646 11935 21042 11936
rect 1761 11658 1827 11661
rect 14457 11658 14523 11661
rect 1761 11656 14523 11658
rect 1761 11600 1766 11656
rect 1822 11600 14462 11656
rect 14518 11600 14523 11656
rect 1761 11598 14523 11600
rect 1761 11595 1827 11598
rect 14457 11595 14523 11598
rect 23197 11658 23263 11661
rect 24200 11658 25000 11688
rect 23197 11656 25000 11658
rect 23197 11600 23202 11656
rect 23258 11600 25000 11656
rect 23197 11598 25000 11600
rect 23197 11595 23263 11598
rect 24200 11568 25000 11598
rect 1906 11456 2302 11457
rect 1906 11392 1912 11456
rect 1976 11392 1992 11456
rect 2056 11392 2072 11456
rect 2136 11392 2152 11456
rect 2216 11392 2232 11456
rect 2296 11392 2302 11456
rect 1906 11391 2302 11392
rect 7906 11456 8302 11457
rect 7906 11392 7912 11456
rect 7976 11392 7992 11456
rect 8056 11392 8072 11456
rect 8136 11392 8152 11456
rect 8216 11392 8232 11456
rect 8296 11392 8302 11456
rect 7906 11391 8302 11392
rect 13906 11456 14302 11457
rect 13906 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14152 11456
rect 14216 11392 14232 11456
rect 14296 11392 14302 11456
rect 13906 11391 14302 11392
rect 19906 11456 20302 11457
rect 19906 11392 19912 11456
rect 19976 11392 19992 11456
rect 20056 11392 20072 11456
rect 20136 11392 20152 11456
rect 20216 11392 20232 11456
rect 20296 11392 20302 11456
rect 19906 11391 20302 11392
rect 21081 11250 21147 11253
rect 23105 11250 23171 11253
rect 21081 11248 23171 11250
rect 21081 11192 21086 11248
rect 21142 11192 23110 11248
rect 23166 11192 23171 11248
rect 21081 11190 23171 11192
rect 21081 11187 21147 11190
rect 23105 11187 23171 11190
rect 0 10978 800 11008
rect 22461 10978 22527 10981
rect 24200 10978 25000 11008
rect 0 10918 1410 10978
rect 0 10888 800 10918
rect 1350 10706 1410 10918
rect 22461 10976 25000 10978
rect 22461 10920 22466 10976
rect 22522 10920 25000 10976
rect 22461 10918 25000 10920
rect 22461 10915 22527 10918
rect 2646 10912 3042 10913
rect 2646 10848 2652 10912
rect 2716 10848 2732 10912
rect 2796 10848 2812 10912
rect 2876 10848 2892 10912
rect 2956 10848 2972 10912
rect 3036 10848 3042 10912
rect 2646 10847 3042 10848
rect 8646 10912 9042 10913
rect 8646 10848 8652 10912
rect 8716 10848 8732 10912
rect 8796 10848 8812 10912
rect 8876 10848 8892 10912
rect 8956 10848 8972 10912
rect 9036 10848 9042 10912
rect 8646 10847 9042 10848
rect 14646 10912 15042 10913
rect 14646 10848 14652 10912
rect 14716 10848 14732 10912
rect 14796 10848 14812 10912
rect 14876 10848 14892 10912
rect 14956 10848 14972 10912
rect 15036 10848 15042 10912
rect 14646 10847 15042 10848
rect 20646 10912 21042 10913
rect 20646 10848 20652 10912
rect 20716 10848 20732 10912
rect 20796 10848 20812 10912
rect 20876 10848 20892 10912
rect 20956 10848 20972 10912
rect 21036 10848 21042 10912
rect 24200 10888 25000 10918
rect 20646 10847 21042 10848
rect 4797 10706 4863 10709
rect 1350 10704 4863 10706
rect 1350 10648 4802 10704
rect 4858 10648 4863 10704
rect 1350 10646 4863 10648
rect 4797 10643 4863 10646
rect 9305 10706 9371 10709
rect 9438 10706 9444 10708
rect 9305 10704 9444 10706
rect 9305 10648 9310 10704
rect 9366 10648 9444 10704
rect 9305 10646 9444 10648
rect 9305 10643 9371 10646
rect 9438 10644 9444 10646
rect 9508 10644 9514 10708
rect 19793 10570 19859 10573
rect 22737 10570 22803 10573
rect 19793 10568 22803 10570
rect 19793 10512 19798 10568
rect 19854 10512 22742 10568
rect 22798 10512 22803 10568
rect 19793 10510 22803 10512
rect 19793 10507 19859 10510
rect 22737 10507 22803 10510
rect 1906 10368 2302 10369
rect 1906 10304 1912 10368
rect 1976 10304 1992 10368
rect 2056 10304 2072 10368
rect 2136 10304 2152 10368
rect 2216 10304 2232 10368
rect 2296 10304 2302 10368
rect 1906 10303 2302 10304
rect 7906 10368 8302 10369
rect 7906 10304 7912 10368
rect 7976 10304 7992 10368
rect 8056 10304 8072 10368
rect 8136 10304 8152 10368
rect 8216 10304 8232 10368
rect 8296 10304 8302 10368
rect 7906 10303 8302 10304
rect 13906 10368 14302 10369
rect 13906 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14152 10368
rect 14216 10304 14232 10368
rect 14296 10304 14302 10368
rect 13906 10303 14302 10304
rect 19906 10368 20302 10369
rect 19906 10304 19912 10368
rect 19976 10304 19992 10368
rect 20056 10304 20072 10368
rect 20136 10304 20152 10368
rect 20216 10304 20232 10368
rect 20296 10304 20302 10368
rect 19906 10303 20302 10304
rect 21173 10298 21239 10301
rect 21449 10298 21515 10301
rect 21173 10296 21515 10298
rect 21173 10240 21178 10296
rect 21234 10240 21454 10296
rect 21510 10240 21515 10296
rect 21173 10238 21515 10240
rect 21173 10235 21239 10238
rect 21449 10235 21515 10238
rect 21265 10162 21331 10165
rect 22277 10162 22343 10165
rect 21265 10160 22343 10162
rect 21265 10104 21270 10160
rect 21326 10104 22282 10160
rect 22338 10104 22343 10160
rect 21265 10102 22343 10104
rect 21265 10099 21331 10102
rect 22277 10099 22343 10102
rect 12617 10026 12683 10029
rect 15469 10026 15535 10029
rect 12617 10024 15535 10026
rect 12617 9968 12622 10024
rect 12678 9968 15474 10024
rect 15530 9968 15535 10024
rect 12617 9966 15535 9968
rect 12617 9963 12683 9966
rect 15469 9963 15535 9966
rect 2646 9824 3042 9825
rect 2646 9760 2652 9824
rect 2716 9760 2732 9824
rect 2796 9760 2812 9824
rect 2876 9760 2892 9824
rect 2956 9760 2972 9824
rect 3036 9760 3042 9824
rect 2646 9759 3042 9760
rect 8646 9824 9042 9825
rect 8646 9760 8652 9824
rect 8716 9760 8732 9824
rect 8796 9760 8812 9824
rect 8876 9760 8892 9824
rect 8956 9760 8972 9824
rect 9036 9760 9042 9824
rect 8646 9759 9042 9760
rect 14646 9824 15042 9825
rect 14646 9760 14652 9824
rect 14716 9760 14732 9824
rect 14796 9760 14812 9824
rect 14876 9760 14892 9824
rect 14956 9760 14972 9824
rect 15036 9760 15042 9824
rect 14646 9759 15042 9760
rect 20646 9824 21042 9825
rect 20646 9760 20652 9824
rect 20716 9760 20732 9824
rect 20796 9760 20812 9824
rect 20876 9760 20892 9824
rect 20956 9760 20972 9824
rect 21036 9760 21042 9824
rect 20646 9759 21042 9760
rect 2221 9618 2287 9621
rect 6453 9618 6519 9621
rect 2221 9616 6519 9618
rect 2221 9560 2226 9616
rect 2282 9560 6458 9616
rect 6514 9560 6519 9616
rect 2221 9558 6519 9560
rect 2221 9555 2287 9558
rect 6453 9555 6519 9558
rect 11237 9618 11303 9621
rect 11881 9618 11947 9621
rect 11237 9616 11947 9618
rect 11237 9560 11242 9616
rect 11298 9560 11886 9616
rect 11942 9560 11947 9616
rect 11237 9558 11947 9560
rect 11237 9555 11303 9558
rect 11881 9555 11947 9558
rect 20805 9618 20871 9621
rect 21173 9618 21239 9621
rect 21725 9618 21791 9621
rect 20805 9616 21239 9618
rect 20805 9560 20810 9616
rect 20866 9560 21178 9616
rect 21234 9560 21239 9616
rect 20805 9558 21239 9560
rect 20805 9555 20871 9558
rect 21173 9555 21239 9558
rect 21406 9616 21791 9618
rect 21406 9560 21730 9616
rect 21786 9560 21791 9616
rect 21406 9558 21791 9560
rect 21406 9485 21466 9558
rect 21725 9555 21791 9558
rect 2405 9482 2471 9485
rect 12433 9482 12499 9485
rect 2405 9480 12499 9482
rect 2405 9424 2410 9480
rect 2466 9424 12438 9480
rect 12494 9424 12499 9480
rect 2405 9422 12499 9424
rect 2405 9419 2471 9422
rect 12433 9419 12499 9422
rect 20069 9482 20135 9485
rect 21357 9482 21466 9485
rect 20069 9480 21466 9482
rect 20069 9424 20074 9480
rect 20130 9424 21362 9480
rect 21418 9424 21466 9480
rect 20069 9422 21466 9424
rect 21633 9482 21699 9485
rect 23289 9482 23355 9485
rect 21633 9480 23355 9482
rect 21633 9424 21638 9480
rect 21694 9424 23294 9480
rect 23350 9424 23355 9480
rect 21633 9422 23355 9424
rect 20069 9419 20135 9422
rect 21357 9419 21423 9422
rect 21633 9419 21699 9422
rect 23289 9419 23355 9422
rect 1906 9280 2302 9281
rect 1906 9216 1912 9280
rect 1976 9216 1992 9280
rect 2056 9216 2072 9280
rect 2136 9216 2152 9280
rect 2216 9216 2232 9280
rect 2296 9216 2302 9280
rect 1906 9215 2302 9216
rect 7906 9280 8302 9281
rect 7906 9216 7912 9280
rect 7976 9216 7992 9280
rect 8056 9216 8072 9280
rect 8136 9216 8152 9280
rect 8216 9216 8232 9280
rect 8296 9216 8302 9280
rect 7906 9215 8302 9216
rect 13906 9280 14302 9281
rect 13906 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14152 9280
rect 14216 9216 14232 9280
rect 14296 9216 14302 9280
rect 13906 9215 14302 9216
rect 19906 9280 20302 9281
rect 19906 9216 19912 9280
rect 19976 9216 19992 9280
rect 20056 9216 20072 9280
rect 20136 9216 20152 9280
rect 20216 9216 20232 9280
rect 20296 9216 20302 9280
rect 19906 9215 20302 9216
rect 23013 8938 23079 8941
rect 24200 8938 25000 8968
rect 23013 8936 25000 8938
rect 23013 8880 23018 8936
rect 23074 8880 25000 8936
rect 23013 8878 25000 8880
rect 23013 8875 23079 8878
rect 24200 8848 25000 8878
rect 2646 8736 3042 8737
rect 2646 8672 2652 8736
rect 2716 8672 2732 8736
rect 2796 8672 2812 8736
rect 2876 8672 2892 8736
rect 2956 8672 2972 8736
rect 3036 8672 3042 8736
rect 2646 8671 3042 8672
rect 8646 8736 9042 8737
rect 8646 8672 8652 8736
rect 8716 8672 8732 8736
rect 8796 8672 8812 8736
rect 8876 8672 8892 8736
rect 8956 8672 8972 8736
rect 9036 8672 9042 8736
rect 8646 8671 9042 8672
rect 14646 8736 15042 8737
rect 14646 8672 14652 8736
rect 14716 8672 14732 8736
rect 14796 8672 14812 8736
rect 14876 8672 14892 8736
rect 14956 8672 14972 8736
rect 15036 8672 15042 8736
rect 14646 8671 15042 8672
rect 20646 8736 21042 8737
rect 20646 8672 20652 8736
rect 20716 8672 20732 8736
rect 20796 8672 20812 8736
rect 20876 8672 20892 8736
rect 20956 8672 20972 8736
rect 21036 8672 21042 8736
rect 20646 8671 21042 8672
rect 23289 8258 23355 8261
rect 24200 8258 25000 8288
rect 23289 8256 25000 8258
rect 23289 8200 23294 8256
rect 23350 8200 25000 8256
rect 23289 8198 25000 8200
rect 23289 8195 23355 8198
rect 1906 8192 2302 8193
rect 1906 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2302 8192
rect 1906 8127 2302 8128
rect 7906 8192 8302 8193
rect 7906 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8072 8192
rect 8136 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8302 8192
rect 7906 8127 8302 8128
rect 13906 8192 14302 8193
rect 13906 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14152 8192
rect 14216 8128 14232 8192
rect 14296 8128 14302 8192
rect 13906 8127 14302 8128
rect 19906 8192 20302 8193
rect 19906 8128 19912 8192
rect 19976 8128 19992 8192
rect 20056 8128 20072 8192
rect 20136 8128 20152 8192
rect 20216 8128 20232 8192
rect 20296 8128 20302 8192
rect 24200 8168 25000 8198
rect 19906 8127 20302 8128
rect 1209 7986 1275 7989
rect 2589 7986 2655 7989
rect 1209 7984 2655 7986
rect 1209 7928 1214 7984
rect 1270 7928 2594 7984
rect 2650 7928 2655 7984
rect 1209 7926 2655 7928
rect 1209 7923 1275 7926
rect 2589 7923 2655 7926
rect 7097 7986 7163 7989
rect 12157 7986 12223 7989
rect 7097 7984 12223 7986
rect 7097 7928 7102 7984
rect 7158 7928 12162 7984
rect 12218 7928 12223 7984
rect 7097 7926 12223 7928
rect 7097 7923 7163 7926
rect 12157 7923 12223 7926
rect 1669 7850 1735 7853
rect 8569 7850 8635 7853
rect 1669 7848 8635 7850
rect 1669 7792 1674 7848
rect 1730 7792 8574 7848
rect 8630 7792 8635 7848
rect 1669 7790 8635 7792
rect 1669 7787 1735 7790
rect 8569 7787 8635 7790
rect 3785 7714 3851 7717
rect 4797 7714 4863 7717
rect 3785 7712 4863 7714
rect 3785 7656 3790 7712
rect 3846 7656 4802 7712
rect 4858 7656 4863 7712
rect 3785 7654 4863 7656
rect 3785 7651 3851 7654
rect 4797 7651 4863 7654
rect 2646 7648 3042 7649
rect 2646 7584 2652 7648
rect 2716 7584 2732 7648
rect 2796 7584 2812 7648
rect 2876 7584 2892 7648
rect 2956 7584 2972 7648
rect 3036 7584 3042 7648
rect 2646 7583 3042 7584
rect 8646 7648 9042 7649
rect 8646 7584 8652 7648
rect 8716 7584 8732 7648
rect 8796 7584 8812 7648
rect 8876 7584 8892 7648
rect 8956 7584 8972 7648
rect 9036 7584 9042 7648
rect 8646 7583 9042 7584
rect 14646 7648 15042 7649
rect 14646 7584 14652 7648
rect 14716 7584 14732 7648
rect 14796 7584 14812 7648
rect 14876 7584 14892 7648
rect 14956 7584 14972 7648
rect 15036 7584 15042 7648
rect 14646 7583 15042 7584
rect 20646 7648 21042 7649
rect 20646 7584 20652 7648
rect 20716 7584 20732 7648
rect 20796 7584 20812 7648
rect 20876 7584 20892 7648
rect 20956 7584 20972 7648
rect 21036 7584 21042 7648
rect 20646 7583 21042 7584
rect 3049 7306 3115 7309
rect 4337 7306 4403 7309
rect 3049 7304 4403 7306
rect 3049 7248 3054 7304
rect 3110 7248 4342 7304
rect 4398 7248 4403 7304
rect 3049 7246 4403 7248
rect 3049 7243 3115 7246
rect 4337 7243 4403 7246
rect 2681 7170 2747 7173
rect 5441 7170 5507 7173
rect 2681 7168 5507 7170
rect 2681 7112 2686 7168
rect 2742 7112 5446 7168
rect 5502 7112 5507 7168
rect 2681 7110 5507 7112
rect 2681 7107 2747 7110
rect 5441 7107 5507 7110
rect 1906 7104 2302 7105
rect 1906 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2302 7104
rect 1906 7039 2302 7040
rect 7906 7104 8302 7105
rect 7906 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8072 7104
rect 8136 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8302 7104
rect 7906 7039 8302 7040
rect 13906 7104 14302 7105
rect 13906 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14152 7104
rect 14216 7040 14232 7104
rect 14296 7040 14302 7104
rect 13906 7039 14302 7040
rect 19906 7104 20302 7105
rect 19906 7040 19912 7104
rect 19976 7040 19992 7104
rect 20056 7040 20072 7104
rect 20136 7040 20152 7104
rect 20216 7040 20232 7104
rect 20296 7040 20302 7104
rect 19906 7039 20302 7040
rect 2773 7034 2839 7037
rect 5349 7034 5415 7037
rect 2773 7032 5415 7034
rect 2773 6976 2778 7032
rect 2834 6976 5354 7032
rect 5410 6976 5415 7032
rect 2773 6974 5415 6976
rect 2773 6971 2839 6974
rect 5349 6971 5415 6974
rect 3049 6898 3115 6901
rect 4521 6898 4587 6901
rect 3049 6896 4587 6898
rect 3049 6840 3054 6896
rect 3110 6840 4526 6896
rect 4582 6840 4587 6896
rect 3049 6838 4587 6840
rect 3049 6835 3115 6838
rect 4521 6835 4587 6838
rect 4613 6762 4679 6765
rect 7005 6762 7071 6765
rect 11237 6762 11303 6765
rect 4613 6760 7071 6762
rect 4613 6704 4618 6760
rect 4674 6704 7010 6760
rect 7066 6704 7071 6760
rect 4613 6702 7071 6704
rect 4613 6699 4679 6702
rect 7005 6699 7071 6702
rect 7238 6760 11303 6762
rect 7238 6704 11242 6760
rect 11298 6704 11303 6760
rect 7238 6702 11303 6704
rect 3969 6626 4035 6629
rect 7238 6626 7298 6702
rect 11237 6699 11303 6702
rect 3969 6624 7298 6626
rect 3969 6568 3974 6624
rect 4030 6568 7298 6624
rect 3969 6566 7298 6568
rect 3969 6563 4035 6566
rect 2646 6560 3042 6561
rect 2646 6496 2652 6560
rect 2716 6496 2732 6560
rect 2796 6496 2812 6560
rect 2876 6496 2892 6560
rect 2956 6496 2972 6560
rect 3036 6496 3042 6560
rect 2646 6495 3042 6496
rect 8646 6560 9042 6561
rect 8646 6496 8652 6560
rect 8716 6496 8732 6560
rect 8796 6496 8812 6560
rect 8876 6496 8892 6560
rect 8956 6496 8972 6560
rect 9036 6496 9042 6560
rect 8646 6495 9042 6496
rect 14646 6560 15042 6561
rect 14646 6496 14652 6560
rect 14716 6496 14732 6560
rect 14796 6496 14812 6560
rect 14876 6496 14892 6560
rect 14956 6496 14972 6560
rect 15036 6496 15042 6560
rect 14646 6495 15042 6496
rect 20646 6560 21042 6561
rect 20646 6496 20652 6560
rect 20716 6496 20732 6560
rect 20796 6496 20812 6560
rect 20876 6496 20892 6560
rect 20956 6496 20972 6560
rect 21036 6496 21042 6560
rect 20646 6495 21042 6496
rect 3785 6490 3851 6493
rect 6913 6490 6979 6493
rect 3785 6488 6979 6490
rect 3785 6432 3790 6488
rect 3846 6432 6918 6488
rect 6974 6432 6979 6488
rect 3785 6430 6979 6432
rect 3785 6427 3851 6430
rect 6913 6427 6979 6430
rect 3049 6354 3115 6357
rect 6729 6354 6795 6357
rect 3049 6352 6795 6354
rect 3049 6296 3054 6352
rect 3110 6296 6734 6352
rect 6790 6296 6795 6352
rect 3049 6294 6795 6296
rect 3049 6291 3115 6294
rect 6729 6291 6795 6294
rect 3049 6218 3115 6221
rect 3509 6218 3575 6221
rect 8293 6218 8359 6221
rect 3049 6216 3575 6218
rect 3049 6160 3054 6216
rect 3110 6160 3514 6216
rect 3570 6160 3575 6216
rect 3049 6158 3575 6160
rect 3049 6155 3115 6158
rect 3509 6155 3575 6158
rect 3742 6216 8359 6218
rect 3742 6160 8298 6216
rect 8354 6160 8359 6216
rect 3742 6158 8359 6160
rect 2405 6082 2471 6085
rect 3742 6082 3802 6158
rect 8293 6155 8359 6158
rect 2405 6080 3802 6082
rect 2405 6024 2410 6080
rect 2466 6024 3802 6080
rect 2405 6022 3802 6024
rect 2405 6019 2471 6022
rect 1906 6016 2302 6017
rect 1906 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2302 6016
rect 1906 5951 2302 5952
rect 7906 6016 8302 6017
rect 7906 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8072 6016
rect 8136 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8302 6016
rect 7906 5951 8302 5952
rect 13906 6016 14302 6017
rect 13906 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14152 6016
rect 14216 5952 14232 6016
rect 14296 5952 14302 6016
rect 13906 5951 14302 5952
rect 19906 6016 20302 6017
rect 19906 5952 19912 6016
rect 19976 5952 19992 6016
rect 20056 5952 20072 6016
rect 20136 5952 20152 6016
rect 20216 5952 20232 6016
rect 20296 5952 20302 6016
rect 19906 5951 20302 5952
rect 3049 5946 3115 5949
rect 3969 5946 4035 5949
rect 3049 5944 4035 5946
rect 3049 5888 3054 5944
rect 3110 5888 3974 5944
rect 4030 5888 4035 5944
rect 3049 5886 4035 5888
rect 3049 5883 3115 5886
rect 3969 5883 4035 5886
rect 2221 5810 2287 5813
rect 6453 5810 6519 5813
rect 2221 5808 6519 5810
rect 2221 5752 2226 5808
rect 2282 5752 6458 5808
rect 6514 5752 6519 5808
rect 2221 5750 6519 5752
rect 2221 5747 2287 5750
rect 6453 5747 6519 5750
rect 2865 5674 2931 5677
rect 3601 5674 3667 5677
rect 2865 5672 3667 5674
rect 2865 5616 2870 5672
rect 2926 5616 3606 5672
rect 3662 5616 3667 5672
rect 2865 5614 3667 5616
rect 2865 5611 2931 5614
rect 3601 5611 3667 5614
rect 2646 5472 3042 5473
rect 2646 5408 2652 5472
rect 2716 5408 2732 5472
rect 2796 5408 2812 5472
rect 2876 5408 2892 5472
rect 2956 5408 2972 5472
rect 3036 5408 3042 5472
rect 2646 5407 3042 5408
rect 8646 5472 9042 5473
rect 8646 5408 8652 5472
rect 8716 5408 8732 5472
rect 8796 5408 8812 5472
rect 8876 5408 8892 5472
rect 8956 5408 8972 5472
rect 9036 5408 9042 5472
rect 8646 5407 9042 5408
rect 14646 5472 15042 5473
rect 14646 5408 14652 5472
rect 14716 5408 14732 5472
rect 14796 5408 14812 5472
rect 14876 5408 14892 5472
rect 14956 5408 14972 5472
rect 15036 5408 15042 5472
rect 14646 5407 15042 5408
rect 20646 5472 21042 5473
rect 20646 5408 20652 5472
rect 20716 5408 20732 5472
rect 20796 5408 20812 5472
rect 20876 5408 20892 5472
rect 20956 5408 20972 5472
rect 21036 5408 21042 5472
rect 20646 5407 21042 5408
rect 1906 4928 2302 4929
rect 1906 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2302 4928
rect 1906 4863 2302 4864
rect 7906 4928 8302 4929
rect 7906 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8072 4928
rect 8136 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8302 4928
rect 7906 4863 8302 4864
rect 13906 4928 14302 4929
rect 13906 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14152 4928
rect 14216 4864 14232 4928
rect 14296 4864 14302 4928
rect 13906 4863 14302 4864
rect 19906 4928 20302 4929
rect 19906 4864 19912 4928
rect 19976 4864 19992 4928
rect 20056 4864 20072 4928
rect 20136 4864 20152 4928
rect 20216 4864 20232 4928
rect 20296 4864 20302 4928
rect 19906 4863 20302 4864
rect 2646 4384 3042 4385
rect 2646 4320 2652 4384
rect 2716 4320 2732 4384
rect 2796 4320 2812 4384
rect 2876 4320 2892 4384
rect 2956 4320 2972 4384
rect 3036 4320 3042 4384
rect 2646 4319 3042 4320
rect 8646 4384 9042 4385
rect 8646 4320 8652 4384
rect 8716 4320 8732 4384
rect 8796 4320 8812 4384
rect 8876 4320 8892 4384
rect 8956 4320 8972 4384
rect 9036 4320 9042 4384
rect 8646 4319 9042 4320
rect 14646 4384 15042 4385
rect 14646 4320 14652 4384
rect 14716 4320 14732 4384
rect 14796 4320 14812 4384
rect 14876 4320 14892 4384
rect 14956 4320 14972 4384
rect 15036 4320 15042 4384
rect 14646 4319 15042 4320
rect 20646 4384 21042 4385
rect 20646 4320 20652 4384
rect 20716 4320 20732 4384
rect 20796 4320 20812 4384
rect 20876 4320 20892 4384
rect 20956 4320 20972 4384
rect 21036 4320 21042 4384
rect 20646 4319 21042 4320
rect 1906 3840 2302 3841
rect 1906 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2302 3840
rect 1906 3775 2302 3776
rect 7906 3840 8302 3841
rect 7906 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8072 3840
rect 8136 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8302 3840
rect 7906 3775 8302 3776
rect 13906 3840 14302 3841
rect 13906 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14152 3840
rect 14216 3776 14232 3840
rect 14296 3776 14302 3840
rect 13906 3775 14302 3776
rect 19906 3840 20302 3841
rect 19906 3776 19912 3840
rect 19976 3776 19992 3840
rect 20056 3776 20072 3840
rect 20136 3776 20152 3840
rect 20216 3776 20232 3840
rect 20296 3776 20302 3840
rect 19906 3775 20302 3776
rect 2646 3296 3042 3297
rect 2646 3232 2652 3296
rect 2716 3232 2732 3296
rect 2796 3232 2812 3296
rect 2876 3232 2892 3296
rect 2956 3232 2972 3296
rect 3036 3232 3042 3296
rect 2646 3231 3042 3232
rect 8646 3296 9042 3297
rect 8646 3232 8652 3296
rect 8716 3232 8732 3296
rect 8796 3232 8812 3296
rect 8876 3232 8892 3296
rect 8956 3232 8972 3296
rect 9036 3232 9042 3296
rect 8646 3231 9042 3232
rect 14646 3296 15042 3297
rect 14646 3232 14652 3296
rect 14716 3232 14732 3296
rect 14796 3232 14812 3296
rect 14876 3232 14892 3296
rect 14956 3232 14972 3296
rect 15036 3232 15042 3296
rect 14646 3231 15042 3232
rect 20646 3296 21042 3297
rect 20646 3232 20652 3296
rect 20716 3232 20732 3296
rect 20796 3232 20812 3296
rect 20876 3232 20892 3296
rect 20956 3232 20972 3296
rect 21036 3232 21042 3296
rect 20646 3231 21042 3232
rect 1906 2752 2302 2753
rect 1906 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2302 2752
rect 1906 2687 2302 2688
rect 7906 2752 8302 2753
rect 7906 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8072 2752
rect 8136 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8302 2752
rect 7906 2687 8302 2688
rect 13906 2752 14302 2753
rect 13906 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14152 2752
rect 14216 2688 14232 2752
rect 14296 2688 14302 2752
rect 13906 2687 14302 2688
rect 19906 2752 20302 2753
rect 19906 2688 19912 2752
rect 19976 2688 19992 2752
rect 20056 2688 20072 2752
rect 20136 2688 20152 2752
rect 20216 2688 20232 2752
rect 20296 2688 20302 2752
rect 19906 2687 20302 2688
rect 2646 2208 3042 2209
rect 2646 2144 2652 2208
rect 2716 2144 2732 2208
rect 2796 2144 2812 2208
rect 2876 2144 2892 2208
rect 2956 2144 2972 2208
rect 3036 2144 3042 2208
rect 2646 2143 3042 2144
rect 8646 2208 9042 2209
rect 8646 2144 8652 2208
rect 8716 2144 8732 2208
rect 8796 2144 8812 2208
rect 8876 2144 8892 2208
rect 8956 2144 8972 2208
rect 9036 2144 9042 2208
rect 8646 2143 9042 2144
rect 14646 2208 15042 2209
rect 14646 2144 14652 2208
rect 14716 2144 14732 2208
rect 14796 2144 14812 2208
rect 14876 2144 14892 2208
rect 14956 2144 14972 2208
rect 15036 2144 15042 2208
rect 14646 2143 15042 2144
rect 20646 2208 21042 2209
rect 20646 2144 20652 2208
rect 20716 2144 20732 2208
rect 20796 2144 20812 2208
rect 20876 2144 20892 2208
rect 20956 2144 20972 2208
rect 21036 2144 21042 2208
rect 20646 2143 21042 2144
<< via3 >>
rect 1912 24508 1976 24512
rect 1912 24452 1916 24508
rect 1916 24452 1972 24508
rect 1972 24452 1976 24508
rect 1912 24448 1976 24452
rect 1992 24508 2056 24512
rect 1992 24452 1996 24508
rect 1996 24452 2052 24508
rect 2052 24452 2056 24508
rect 1992 24448 2056 24452
rect 2072 24508 2136 24512
rect 2072 24452 2076 24508
rect 2076 24452 2132 24508
rect 2132 24452 2136 24508
rect 2072 24448 2136 24452
rect 2152 24508 2216 24512
rect 2152 24452 2156 24508
rect 2156 24452 2212 24508
rect 2212 24452 2216 24508
rect 2152 24448 2216 24452
rect 2232 24508 2296 24512
rect 2232 24452 2236 24508
rect 2236 24452 2292 24508
rect 2292 24452 2296 24508
rect 2232 24448 2296 24452
rect 7912 24508 7976 24512
rect 7912 24452 7916 24508
rect 7916 24452 7972 24508
rect 7972 24452 7976 24508
rect 7912 24448 7976 24452
rect 7992 24508 8056 24512
rect 7992 24452 7996 24508
rect 7996 24452 8052 24508
rect 8052 24452 8056 24508
rect 7992 24448 8056 24452
rect 8072 24508 8136 24512
rect 8072 24452 8076 24508
rect 8076 24452 8132 24508
rect 8132 24452 8136 24508
rect 8072 24448 8136 24452
rect 8152 24508 8216 24512
rect 8152 24452 8156 24508
rect 8156 24452 8212 24508
rect 8212 24452 8216 24508
rect 8152 24448 8216 24452
rect 8232 24508 8296 24512
rect 8232 24452 8236 24508
rect 8236 24452 8292 24508
rect 8292 24452 8296 24508
rect 8232 24448 8296 24452
rect 13912 24508 13976 24512
rect 13912 24452 13916 24508
rect 13916 24452 13972 24508
rect 13972 24452 13976 24508
rect 13912 24448 13976 24452
rect 13992 24508 14056 24512
rect 13992 24452 13996 24508
rect 13996 24452 14052 24508
rect 14052 24452 14056 24508
rect 13992 24448 14056 24452
rect 14072 24508 14136 24512
rect 14072 24452 14076 24508
rect 14076 24452 14132 24508
rect 14132 24452 14136 24508
rect 14072 24448 14136 24452
rect 14152 24508 14216 24512
rect 14152 24452 14156 24508
rect 14156 24452 14212 24508
rect 14212 24452 14216 24508
rect 14152 24448 14216 24452
rect 14232 24508 14296 24512
rect 14232 24452 14236 24508
rect 14236 24452 14292 24508
rect 14292 24452 14296 24508
rect 14232 24448 14296 24452
rect 19912 24508 19976 24512
rect 19912 24452 19916 24508
rect 19916 24452 19972 24508
rect 19972 24452 19976 24508
rect 19912 24448 19976 24452
rect 19992 24508 20056 24512
rect 19992 24452 19996 24508
rect 19996 24452 20052 24508
rect 20052 24452 20056 24508
rect 19992 24448 20056 24452
rect 20072 24508 20136 24512
rect 20072 24452 20076 24508
rect 20076 24452 20132 24508
rect 20132 24452 20136 24508
rect 20072 24448 20136 24452
rect 20152 24508 20216 24512
rect 20152 24452 20156 24508
rect 20156 24452 20212 24508
rect 20212 24452 20216 24508
rect 20152 24448 20216 24452
rect 20232 24508 20296 24512
rect 20232 24452 20236 24508
rect 20236 24452 20292 24508
rect 20292 24452 20296 24508
rect 20232 24448 20296 24452
rect 2652 23964 2716 23968
rect 2652 23908 2656 23964
rect 2656 23908 2712 23964
rect 2712 23908 2716 23964
rect 2652 23904 2716 23908
rect 2732 23964 2796 23968
rect 2732 23908 2736 23964
rect 2736 23908 2792 23964
rect 2792 23908 2796 23964
rect 2732 23904 2796 23908
rect 2812 23964 2876 23968
rect 2812 23908 2816 23964
rect 2816 23908 2872 23964
rect 2872 23908 2876 23964
rect 2812 23904 2876 23908
rect 2892 23964 2956 23968
rect 2892 23908 2896 23964
rect 2896 23908 2952 23964
rect 2952 23908 2956 23964
rect 2892 23904 2956 23908
rect 2972 23964 3036 23968
rect 2972 23908 2976 23964
rect 2976 23908 3032 23964
rect 3032 23908 3036 23964
rect 2972 23904 3036 23908
rect 8652 23964 8716 23968
rect 8652 23908 8656 23964
rect 8656 23908 8712 23964
rect 8712 23908 8716 23964
rect 8652 23904 8716 23908
rect 8732 23964 8796 23968
rect 8732 23908 8736 23964
rect 8736 23908 8792 23964
rect 8792 23908 8796 23964
rect 8732 23904 8796 23908
rect 8812 23964 8876 23968
rect 8812 23908 8816 23964
rect 8816 23908 8872 23964
rect 8872 23908 8876 23964
rect 8812 23904 8876 23908
rect 8892 23964 8956 23968
rect 8892 23908 8896 23964
rect 8896 23908 8952 23964
rect 8952 23908 8956 23964
rect 8892 23904 8956 23908
rect 8972 23964 9036 23968
rect 8972 23908 8976 23964
rect 8976 23908 9032 23964
rect 9032 23908 9036 23964
rect 8972 23904 9036 23908
rect 14652 23964 14716 23968
rect 14652 23908 14656 23964
rect 14656 23908 14712 23964
rect 14712 23908 14716 23964
rect 14652 23904 14716 23908
rect 14732 23964 14796 23968
rect 14732 23908 14736 23964
rect 14736 23908 14792 23964
rect 14792 23908 14796 23964
rect 14732 23904 14796 23908
rect 14812 23964 14876 23968
rect 14812 23908 14816 23964
rect 14816 23908 14872 23964
rect 14872 23908 14876 23964
rect 14812 23904 14876 23908
rect 14892 23964 14956 23968
rect 14892 23908 14896 23964
rect 14896 23908 14952 23964
rect 14952 23908 14956 23964
rect 14892 23904 14956 23908
rect 14972 23964 15036 23968
rect 14972 23908 14976 23964
rect 14976 23908 15032 23964
rect 15032 23908 15036 23964
rect 14972 23904 15036 23908
rect 20652 23964 20716 23968
rect 20652 23908 20656 23964
rect 20656 23908 20712 23964
rect 20712 23908 20716 23964
rect 20652 23904 20716 23908
rect 20732 23964 20796 23968
rect 20732 23908 20736 23964
rect 20736 23908 20792 23964
rect 20792 23908 20796 23964
rect 20732 23904 20796 23908
rect 20812 23964 20876 23968
rect 20812 23908 20816 23964
rect 20816 23908 20872 23964
rect 20872 23908 20876 23964
rect 20812 23904 20876 23908
rect 20892 23964 20956 23968
rect 20892 23908 20896 23964
rect 20896 23908 20952 23964
rect 20952 23908 20956 23964
rect 20892 23904 20956 23908
rect 20972 23964 21036 23968
rect 20972 23908 20976 23964
rect 20976 23908 21032 23964
rect 21032 23908 21036 23964
rect 20972 23904 21036 23908
rect 1912 23420 1976 23424
rect 1912 23364 1916 23420
rect 1916 23364 1972 23420
rect 1972 23364 1976 23420
rect 1912 23360 1976 23364
rect 1992 23420 2056 23424
rect 1992 23364 1996 23420
rect 1996 23364 2052 23420
rect 2052 23364 2056 23420
rect 1992 23360 2056 23364
rect 2072 23420 2136 23424
rect 2072 23364 2076 23420
rect 2076 23364 2132 23420
rect 2132 23364 2136 23420
rect 2072 23360 2136 23364
rect 2152 23420 2216 23424
rect 2152 23364 2156 23420
rect 2156 23364 2212 23420
rect 2212 23364 2216 23420
rect 2152 23360 2216 23364
rect 2232 23420 2296 23424
rect 2232 23364 2236 23420
rect 2236 23364 2292 23420
rect 2292 23364 2296 23420
rect 2232 23360 2296 23364
rect 7912 23420 7976 23424
rect 7912 23364 7916 23420
rect 7916 23364 7972 23420
rect 7972 23364 7976 23420
rect 7912 23360 7976 23364
rect 7992 23420 8056 23424
rect 7992 23364 7996 23420
rect 7996 23364 8052 23420
rect 8052 23364 8056 23420
rect 7992 23360 8056 23364
rect 8072 23420 8136 23424
rect 8072 23364 8076 23420
rect 8076 23364 8132 23420
rect 8132 23364 8136 23420
rect 8072 23360 8136 23364
rect 8152 23420 8216 23424
rect 8152 23364 8156 23420
rect 8156 23364 8212 23420
rect 8212 23364 8216 23420
rect 8152 23360 8216 23364
rect 8232 23420 8296 23424
rect 8232 23364 8236 23420
rect 8236 23364 8292 23420
rect 8292 23364 8296 23420
rect 8232 23360 8296 23364
rect 13912 23420 13976 23424
rect 13912 23364 13916 23420
rect 13916 23364 13972 23420
rect 13972 23364 13976 23420
rect 13912 23360 13976 23364
rect 13992 23420 14056 23424
rect 13992 23364 13996 23420
rect 13996 23364 14052 23420
rect 14052 23364 14056 23420
rect 13992 23360 14056 23364
rect 14072 23420 14136 23424
rect 14072 23364 14076 23420
rect 14076 23364 14132 23420
rect 14132 23364 14136 23420
rect 14072 23360 14136 23364
rect 14152 23420 14216 23424
rect 14152 23364 14156 23420
rect 14156 23364 14212 23420
rect 14212 23364 14216 23420
rect 14152 23360 14216 23364
rect 14232 23420 14296 23424
rect 14232 23364 14236 23420
rect 14236 23364 14292 23420
rect 14292 23364 14296 23420
rect 14232 23360 14296 23364
rect 19912 23420 19976 23424
rect 19912 23364 19916 23420
rect 19916 23364 19972 23420
rect 19972 23364 19976 23420
rect 19912 23360 19976 23364
rect 19992 23420 20056 23424
rect 19992 23364 19996 23420
rect 19996 23364 20052 23420
rect 20052 23364 20056 23420
rect 19992 23360 20056 23364
rect 20072 23420 20136 23424
rect 20072 23364 20076 23420
rect 20076 23364 20132 23420
rect 20132 23364 20136 23420
rect 20072 23360 20136 23364
rect 20152 23420 20216 23424
rect 20152 23364 20156 23420
rect 20156 23364 20212 23420
rect 20212 23364 20216 23420
rect 20152 23360 20216 23364
rect 20232 23420 20296 23424
rect 20232 23364 20236 23420
rect 20236 23364 20292 23420
rect 20292 23364 20296 23420
rect 20232 23360 20296 23364
rect 2652 22876 2716 22880
rect 2652 22820 2656 22876
rect 2656 22820 2712 22876
rect 2712 22820 2716 22876
rect 2652 22816 2716 22820
rect 2732 22876 2796 22880
rect 2732 22820 2736 22876
rect 2736 22820 2792 22876
rect 2792 22820 2796 22876
rect 2732 22816 2796 22820
rect 2812 22876 2876 22880
rect 2812 22820 2816 22876
rect 2816 22820 2872 22876
rect 2872 22820 2876 22876
rect 2812 22816 2876 22820
rect 2892 22876 2956 22880
rect 2892 22820 2896 22876
rect 2896 22820 2952 22876
rect 2952 22820 2956 22876
rect 2892 22816 2956 22820
rect 2972 22876 3036 22880
rect 2972 22820 2976 22876
rect 2976 22820 3032 22876
rect 3032 22820 3036 22876
rect 2972 22816 3036 22820
rect 8652 22876 8716 22880
rect 8652 22820 8656 22876
rect 8656 22820 8712 22876
rect 8712 22820 8716 22876
rect 8652 22816 8716 22820
rect 8732 22876 8796 22880
rect 8732 22820 8736 22876
rect 8736 22820 8792 22876
rect 8792 22820 8796 22876
rect 8732 22816 8796 22820
rect 8812 22876 8876 22880
rect 8812 22820 8816 22876
rect 8816 22820 8872 22876
rect 8872 22820 8876 22876
rect 8812 22816 8876 22820
rect 8892 22876 8956 22880
rect 8892 22820 8896 22876
rect 8896 22820 8952 22876
rect 8952 22820 8956 22876
rect 8892 22816 8956 22820
rect 8972 22876 9036 22880
rect 8972 22820 8976 22876
rect 8976 22820 9032 22876
rect 9032 22820 9036 22876
rect 8972 22816 9036 22820
rect 14652 22876 14716 22880
rect 14652 22820 14656 22876
rect 14656 22820 14712 22876
rect 14712 22820 14716 22876
rect 14652 22816 14716 22820
rect 14732 22876 14796 22880
rect 14732 22820 14736 22876
rect 14736 22820 14792 22876
rect 14792 22820 14796 22876
rect 14732 22816 14796 22820
rect 14812 22876 14876 22880
rect 14812 22820 14816 22876
rect 14816 22820 14872 22876
rect 14872 22820 14876 22876
rect 14812 22816 14876 22820
rect 14892 22876 14956 22880
rect 14892 22820 14896 22876
rect 14896 22820 14952 22876
rect 14952 22820 14956 22876
rect 14892 22816 14956 22820
rect 14972 22876 15036 22880
rect 14972 22820 14976 22876
rect 14976 22820 15032 22876
rect 15032 22820 15036 22876
rect 14972 22816 15036 22820
rect 20652 22876 20716 22880
rect 20652 22820 20656 22876
rect 20656 22820 20712 22876
rect 20712 22820 20716 22876
rect 20652 22816 20716 22820
rect 20732 22876 20796 22880
rect 20732 22820 20736 22876
rect 20736 22820 20792 22876
rect 20792 22820 20796 22876
rect 20732 22816 20796 22820
rect 20812 22876 20876 22880
rect 20812 22820 20816 22876
rect 20816 22820 20872 22876
rect 20872 22820 20876 22876
rect 20812 22816 20876 22820
rect 20892 22876 20956 22880
rect 20892 22820 20896 22876
rect 20896 22820 20952 22876
rect 20952 22820 20956 22876
rect 20892 22816 20956 22820
rect 20972 22876 21036 22880
rect 20972 22820 20976 22876
rect 20976 22820 21032 22876
rect 21032 22820 21036 22876
rect 20972 22816 21036 22820
rect 1912 22332 1976 22336
rect 1912 22276 1916 22332
rect 1916 22276 1972 22332
rect 1972 22276 1976 22332
rect 1912 22272 1976 22276
rect 1992 22332 2056 22336
rect 1992 22276 1996 22332
rect 1996 22276 2052 22332
rect 2052 22276 2056 22332
rect 1992 22272 2056 22276
rect 2072 22332 2136 22336
rect 2072 22276 2076 22332
rect 2076 22276 2132 22332
rect 2132 22276 2136 22332
rect 2072 22272 2136 22276
rect 2152 22332 2216 22336
rect 2152 22276 2156 22332
rect 2156 22276 2212 22332
rect 2212 22276 2216 22332
rect 2152 22272 2216 22276
rect 2232 22332 2296 22336
rect 2232 22276 2236 22332
rect 2236 22276 2292 22332
rect 2292 22276 2296 22332
rect 2232 22272 2296 22276
rect 7912 22332 7976 22336
rect 7912 22276 7916 22332
rect 7916 22276 7972 22332
rect 7972 22276 7976 22332
rect 7912 22272 7976 22276
rect 7992 22332 8056 22336
rect 7992 22276 7996 22332
rect 7996 22276 8052 22332
rect 8052 22276 8056 22332
rect 7992 22272 8056 22276
rect 8072 22332 8136 22336
rect 8072 22276 8076 22332
rect 8076 22276 8132 22332
rect 8132 22276 8136 22332
rect 8072 22272 8136 22276
rect 8152 22332 8216 22336
rect 8152 22276 8156 22332
rect 8156 22276 8212 22332
rect 8212 22276 8216 22332
rect 8152 22272 8216 22276
rect 8232 22332 8296 22336
rect 8232 22276 8236 22332
rect 8236 22276 8292 22332
rect 8292 22276 8296 22332
rect 8232 22272 8296 22276
rect 13912 22332 13976 22336
rect 13912 22276 13916 22332
rect 13916 22276 13972 22332
rect 13972 22276 13976 22332
rect 13912 22272 13976 22276
rect 13992 22332 14056 22336
rect 13992 22276 13996 22332
rect 13996 22276 14052 22332
rect 14052 22276 14056 22332
rect 13992 22272 14056 22276
rect 14072 22332 14136 22336
rect 14072 22276 14076 22332
rect 14076 22276 14132 22332
rect 14132 22276 14136 22332
rect 14072 22272 14136 22276
rect 14152 22332 14216 22336
rect 14152 22276 14156 22332
rect 14156 22276 14212 22332
rect 14212 22276 14216 22332
rect 14152 22272 14216 22276
rect 14232 22332 14296 22336
rect 14232 22276 14236 22332
rect 14236 22276 14292 22332
rect 14292 22276 14296 22332
rect 14232 22272 14296 22276
rect 19912 22332 19976 22336
rect 19912 22276 19916 22332
rect 19916 22276 19972 22332
rect 19972 22276 19976 22332
rect 19912 22272 19976 22276
rect 19992 22332 20056 22336
rect 19992 22276 19996 22332
rect 19996 22276 20052 22332
rect 20052 22276 20056 22332
rect 19992 22272 20056 22276
rect 20072 22332 20136 22336
rect 20072 22276 20076 22332
rect 20076 22276 20132 22332
rect 20132 22276 20136 22332
rect 20072 22272 20136 22276
rect 20152 22332 20216 22336
rect 20152 22276 20156 22332
rect 20156 22276 20212 22332
rect 20212 22276 20216 22332
rect 20152 22272 20216 22276
rect 20232 22332 20296 22336
rect 20232 22276 20236 22332
rect 20236 22276 20292 22332
rect 20292 22276 20296 22332
rect 20232 22272 20296 22276
rect 2652 21788 2716 21792
rect 2652 21732 2656 21788
rect 2656 21732 2712 21788
rect 2712 21732 2716 21788
rect 2652 21728 2716 21732
rect 2732 21788 2796 21792
rect 2732 21732 2736 21788
rect 2736 21732 2792 21788
rect 2792 21732 2796 21788
rect 2732 21728 2796 21732
rect 2812 21788 2876 21792
rect 2812 21732 2816 21788
rect 2816 21732 2872 21788
rect 2872 21732 2876 21788
rect 2812 21728 2876 21732
rect 2892 21788 2956 21792
rect 2892 21732 2896 21788
rect 2896 21732 2952 21788
rect 2952 21732 2956 21788
rect 2892 21728 2956 21732
rect 2972 21788 3036 21792
rect 2972 21732 2976 21788
rect 2976 21732 3032 21788
rect 3032 21732 3036 21788
rect 2972 21728 3036 21732
rect 8652 21788 8716 21792
rect 8652 21732 8656 21788
rect 8656 21732 8712 21788
rect 8712 21732 8716 21788
rect 8652 21728 8716 21732
rect 8732 21788 8796 21792
rect 8732 21732 8736 21788
rect 8736 21732 8792 21788
rect 8792 21732 8796 21788
rect 8732 21728 8796 21732
rect 8812 21788 8876 21792
rect 8812 21732 8816 21788
rect 8816 21732 8872 21788
rect 8872 21732 8876 21788
rect 8812 21728 8876 21732
rect 8892 21788 8956 21792
rect 8892 21732 8896 21788
rect 8896 21732 8952 21788
rect 8952 21732 8956 21788
rect 8892 21728 8956 21732
rect 8972 21788 9036 21792
rect 8972 21732 8976 21788
rect 8976 21732 9032 21788
rect 9032 21732 9036 21788
rect 8972 21728 9036 21732
rect 14652 21788 14716 21792
rect 14652 21732 14656 21788
rect 14656 21732 14712 21788
rect 14712 21732 14716 21788
rect 14652 21728 14716 21732
rect 14732 21788 14796 21792
rect 14732 21732 14736 21788
rect 14736 21732 14792 21788
rect 14792 21732 14796 21788
rect 14732 21728 14796 21732
rect 14812 21788 14876 21792
rect 14812 21732 14816 21788
rect 14816 21732 14872 21788
rect 14872 21732 14876 21788
rect 14812 21728 14876 21732
rect 14892 21788 14956 21792
rect 14892 21732 14896 21788
rect 14896 21732 14952 21788
rect 14952 21732 14956 21788
rect 14892 21728 14956 21732
rect 14972 21788 15036 21792
rect 14972 21732 14976 21788
rect 14976 21732 15032 21788
rect 15032 21732 15036 21788
rect 14972 21728 15036 21732
rect 20652 21788 20716 21792
rect 20652 21732 20656 21788
rect 20656 21732 20712 21788
rect 20712 21732 20716 21788
rect 20652 21728 20716 21732
rect 20732 21788 20796 21792
rect 20732 21732 20736 21788
rect 20736 21732 20792 21788
rect 20792 21732 20796 21788
rect 20732 21728 20796 21732
rect 20812 21788 20876 21792
rect 20812 21732 20816 21788
rect 20816 21732 20872 21788
rect 20872 21732 20876 21788
rect 20812 21728 20876 21732
rect 20892 21788 20956 21792
rect 20892 21732 20896 21788
rect 20896 21732 20952 21788
rect 20952 21732 20956 21788
rect 20892 21728 20956 21732
rect 20972 21788 21036 21792
rect 20972 21732 20976 21788
rect 20976 21732 21032 21788
rect 21032 21732 21036 21788
rect 20972 21728 21036 21732
rect 1912 21244 1976 21248
rect 1912 21188 1916 21244
rect 1916 21188 1972 21244
rect 1972 21188 1976 21244
rect 1912 21184 1976 21188
rect 1992 21244 2056 21248
rect 1992 21188 1996 21244
rect 1996 21188 2052 21244
rect 2052 21188 2056 21244
rect 1992 21184 2056 21188
rect 2072 21244 2136 21248
rect 2072 21188 2076 21244
rect 2076 21188 2132 21244
rect 2132 21188 2136 21244
rect 2072 21184 2136 21188
rect 2152 21244 2216 21248
rect 2152 21188 2156 21244
rect 2156 21188 2212 21244
rect 2212 21188 2216 21244
rect 2152 21184 2216 21188
rect 2232 21244 2296 21248
rect 2232 21188 2236 21244
rect 2236 21188 2292 21244
rect 2292 21188 2296 21244
rect 2232 21184 2296 21188
rect 7912 21244 7976 21248
rect 7912 21188 7916 21244
rect 7916 21188 7972 21244
rect 7972 21188 7976 21244
rect 7912 21184 7976 21188
rect 7992 21244 8056 21248
rect 7992 21188 7996 21244
rect 7996 21188 8052 21244
rect 8052 21188 8056 21244
rect 7992 21184 8056 21188
rect 8072 21244 8136 21248
rect 8072 21188 8076 21244
rect 8076 21188 8132 21244
rect 8132 21188 8136 21244
rect 8072 21184 8136 21188
rect 8152 21244 8216 21248
rect 8152 21188 8156 21244
rect 8156 21188 8212 21244
rect 8212 21188 8216 21244
rect 8152 21184 8216 21188
rect 8232 21244 8296 21248
rect 8232 21188 8236 21244
rect 8236 21188 8292 21244
rect 8292 21188 8296 21244
rect 8232 21184 8296 21188
rect 13912 21244 13976 21248
rect 13912 21188 13916 21244
rect 13916 21188 13972 21244
rect 13972 21188 13976 21244
rect 13912 21184 13976 21188
rect 13992 21244 14056 21248
rect 13992 21188 13996 21244
rect 13996 21188 14052 21244
rect 14052 21188 14056 21244
rect 13992 21184 14056 21188
rect 14072 21244 14136 21248
rect 14072 21188 14076 21244
rect 14076 21188 14132 21244
rect 14132 21188 14136 21244
rect 14072 21184 14136 21188
rect 14152 21244 14216 21248
rect 14152 21188 14156 21244
rect 14156 21188 14212 21244
rect 14212 21188 14216 21244
rect 14152 21184 14216 21188
rect 14232 21244 14296 21248
rect 14232 21188 14236 21244
rect 14236 21188 14292 21244
rect 14292 21188 14296 21244
rect 14232 21184 14296 21188
rect 19912 21244 19976 21248
rect 19912 21188 19916 21244
rect 19916 21188 19972 21244
rect 19972 21188 19976 21244
rect 19912 21184 19976 21188
rect 19992 21244 20056 21248
rect 19992 21188 19996 21244
rect 19996 21188 20052 21244
rect 20052 21188 20056 21244
rect 19992 21184 20056 21188
rect 20072 21244 20136 21248
rect 20072 21188 20076 21244
rect 20076 21188 20132 21244
rect 20132 21188 20136 21244
rect 20072 21184 20136 21188
rect 20152 21244 20216 21248
rect 20152 21188 20156 21244
rect 20156 21188 20212 21244
rect 20212 21188 20216 21244
rect 20152 21184 20216 21188
rect 20232 21244 20296 21248
rect 20232 21188 20236 21244
rect 20236 21188 20292 21244
rect 20292 21188 20296 21244
rect 20232 21184 20296 21188
rect 2652 20700 2716 20704
rect 2652 20644 2656 20700
rect 2656 20644 2712 20700
rect 2712 20644 2716 20700
rect 2652 20640 2716 20644
rect 2732 20700 2796 20704
rect 2732 20644 2736 20700
rect 2736 20644 2792 20700
rect 2792 20644 2796 20700
rect 2732 20640 2796 20644
rect 2812 20700 2876 20704
rect 2812 20644 2816 20700
rect 2816 20644 2872 20700
rect 2872 20644 2876 20700
rect 2812 20640 2876 20644
rect 2892 20700 2956 20704
rect 2892 20644 2896 20700
rect 2896 20644 2952 20700
rect 2952 20644 2956 20700
rect 2892 20640 2956 20644
rect 2972 20700 3036 20704
rect 2972 20644 2976 20700
rect 2976 20644 3032 20700
rect 3032 20644 3036 20700
rect 2972 20640 3036 20644
rect 8652 20700 8716 20704
rect 8652 20644 8656 20700
rect 8656 20644 8712 20700
rect 8712 20644 8716 20700
rect 8652 20640 8716 20644
rect 8732 20700 8796 20704
rect 8732 20644 8736 20700
rect 8736 20644 8792 20700
rect 8792 20644 8796 20700
rect 8732 20640 8796 20644
rect 8812 20700 8876 20704
rect 8812 20644 8816 20700
rect 8816 20644 8872 20700
rect 8872 20644 8876 20700
rect 8812 20640 8876 20644
rect 8892 20700 8956 20704
rect 8892 20644 8896 20700
rect 8896 20644 8952 20700
rect 8952 20644 8956 20700
rect 8892 20640 8956 20644
rect 8972 20700 9036 20704
rect 8972 20644 8976 20700
rect 8976 20644 9032 20700
rect 9032 20644 9036 20700
rect 8972 20640 9036 20644
rect 14652 20700 14716 20704
rect 14652 20644 14656 20700
rect 14656 20644 14712 20700
rect 14712 20644 14716 20700
rect 14652 20640 14716 20644
rect 14732 20700 14796 20704
rect 14732 20644 14736 20700
rect 14736 20644 14792 20700
rect 14792 20644 14796 20700
rect 14732 20640 14796 20644
rect 14812 20700 14876 20704
rect 14812 20644 14816 20700
rect 14816 20644 14872 20700
rect 14872 20644 14876 20700
rect 14812 20640 14876 20644
rect 14892 20700 14956 20704
rect 14892 20644 14896 20700
rect 14896 20644 14952 20700
rect 14952 20644 14956 20700
rect 14892 20640 14956 20644
rect 14972 20700 15036 20704
rect 14972 20644 14976 20700
rect 14976 20644 15032 20700
rect 15032 20644 15036 20700
rect 14972 20640 15036 20644
rect 20652 20700 20716 20704
rect 20652 20644 20656 20700
rect 20656 20644 20712 20700
rect 20712 20644 20716 20700
rect 20652 20640 20716 20644
rect 20732 20700 20796 20704
rect 20732 20644 20736 20700
rect 20736 20644 20792 20700
rect 20792 20644 20796 20700
rect 20732 20640 20796 20644
rect 20812 20700 20876 20704
rect 20812 20644 20816 20700
rect 20816 20644 20872 20700
rect 20872 20644 20876 20700
rect 20812 20640 20876 20644
rect 20892 20700 20956 20704
rect 20892 20644 20896 20700
rect 20896 20644 20952 20700
rect 20952 20644 20956 20700
rect 20892 20640 20956 20644
rect 20972 20700 21036 20704
rect 20972 20644 20976 20700
rect 20976 20644 21032 20700
rect 21032 20644 21036 20700
rect 20972 20640 21036 20644
rect 1912 20156 1976 20160
rect 1912 20100 1916 20156
rect 1916 20100 1972 20156
rect 1972 20100 1976 20156
rect 1912 20096 1976 20100
rect 1992 20156 2056 20160
rect 1992 20100 1996 20156
rect 1996 20100 2052 20156
rect 2052 20100 2056 20156
rect 1992 20096 2056 20100
rect 2072 20156 2136 20160
rect 2072 20100 2076 20156
rect 2076 20100 2132 20156
rect 2132 20100 2136 20156
rect 2072 20096 2136 20100
rect 2152 20156 2216 20160
rect 2152 20100 2156 20156
rect 2156 20100 2212 20156
rect 2212 20100 2216 20156
rect 2152 20096 2216 20100
rect 2232 20156 2296 20160
rect 2232 20100 2236 20156
rect 2236 20100 2292 20156
rect 2292 20100 2296 20156
rect 2232 20096 2296 20100
rect 7912 20156 7976 20160
rect 7912 20100 7916 20156
rect 7916 20100 7972 20156
rect 7972 20100 7976 20156
rect 7912 20096 7976 20100
rect 7992 20156 8056 20160
rect 7992 20100 7996 20156
rect 7996 20100 8052 20156
rect 8052 20100 8056 20156
rect 7992 20096 8056 20100
rect 8072 20156 8136 20160
rect 8072 20100 8076 20156
rect 8076 20100 8132 20156
rect 8132 20100 8136 20156
rect 8072 20096 8136 20100
rect 8152 20156 8216 20160
rect 8152 20100 8156 20156
rect 8156 20100 8212 20156
rect 8212 20100 8216 20156
rect 8152 20096 8216 20100
rect 8232 20156 8296 20160
rect 8232 20100 8236 20156
rect 8236 20100 8292 20156
rect 8292 20100 8296 20156
rect 8232 20096 8296 20100
rect 13912 20156 13976 20160
rect 13912 20100 13916 20156
rect 13916 20100 13972 20156
rect 13972 20100 13976 20156
rect 13912 20096 13976 20100
rect 13992 20156 14056 20160
rect 13992 20100 13996 20156
rect 13996 20100 14052 20156
rect 14052 20100 14056 20156
rect 13992 20096 14056 20100
rect 14072 20156 14136 20160
rect 14072 20100 14076 20156
rect 14076 20100 14132 20156
rect 14132 20100 14136 20156
rect 14072 20096 14136 20100
rect 14152 20156 14216 20160
rect 14152 20100 14156 20156
rect 14156 20100 14212 20156
rect 14212 20100 14216 20156
rect 14152 20096 14216 20100
rect 14232 20156 14296 20160
rect 14232 20100 14236 20156
rect 14236 20100 14292 20156
rect 14292 20100 14296 20156
rect 14232 20096 14296 20100
rect 19912 20156 19976 20160
rect 19912 20100 19916 20156
rect 19916 20100 19972 20156
rect 19972 20100 19976 20156
rect 19912 20096 19976 20100
rect 19992 20156 20056 20160
rect 19992 20100 19996 20156
rect 19996 20100 20052 20156
rect 20052 20100 20056 20156
rect 19992 20096 20056 20100
rect 20072 20156 20136 20160
rect 20072 20100 20076 20156
rect 20076 20100 20132 20156
rect 20132 20100 20136 20156
rect 20072 20096 20136 20100
rect 20152 20156 20216 20160
rect 20152 20100 20156 20156
rect 20156 20100 20212 20156
rect 20212 20100 20216 20156
rect 20152 20096 20216 20100
rect 20232 20156 20296 20160
rect 20232 20100 20236 20156
rect 20236 20100 20292 20156
rect 20292 20100 20296 20156
rect 20232 20096 20296 20100
rect 2652 19612 2716 19616
rect 2652 19556 2656 19612
rect 2656 19556 2712 19612
rect 2712 19556 2716 19612
rect 2652 19552 2716 19556
rect 2732 19612 2796 19616
rect 2732 19556 2736 19612
rect 2736 19556 2792 19612
rect 2792 19556 2796 19612
rect 2732 19552 2796 19556
rect 2812 19612 2876 19616
rect 2812 19556 2816 19612
rect 2816 19556 2872 19612
rect 2872 19556 2876 19612
rect 2812 19552 2876 19556
rect 2892 19612 2956 19616
rect 2892 19556 2896 19612
rect 2896 19556 2952 19612
rect 2952 19556 2956 19612
rect 2892 19552 2956 19556
rect 2972 19612 3036 19616
rect 2972 19556 2976 19612
rect 2976 19556 3032 19612
rect 3032 19556 3036 19612
rect 2972 19552 3036 19556
rect 8652 19612 8716 19616
rect 8652 19556 8656 19612
rect 8656 19556 8712 19612
rect 8712 19556 8716 19612
rect 8652 19552 8716 19556
rect 8732 19612 8796 19616
rect 8732 19556 8736 19612
rect 8736 19556 8792 19612
rect 8792 19556 8796 19612
rect 8732 19552 8796 19556
rect 8812 19612 8876 19616
rect 8812 19556 8816 19612
rect 8816 19556 8872 19612
rect 8872 19556 8876 19612
rect 8812 19552 8876 19556
rect 8892 19612 8956 19616
rect 8892 19556 8896 19612
rect 8896 19556 8952 19612
rect 8952 19556 8956 19612
rect 8892 19552 8956 19556
rect 8972 19612 9036 19616
rect 8972 19556 8976 19612
rect 8976 19556 9032 19612
rect 9032 19556 9036 19612
rect 8972 19552 9036 19556
rect 14652 19612 14716 19616
rect 14652 19556 14656 19612
rect 14656 19556 14712 19612
rect 14712 19556 14716 19612
rect 14652 19552 14716 19556
rect 14732 19612 14796 19616
rect 14732 19556 14736 19612
rect 14736 19556 14792 19612
rect 14792 19556 14796 19612
rect 14732 19552 14796 19556
rect 14812 19612 14876 19616
rect 14812 19556 14816 19612
rect 14816 19556 14872 19612
rect 14872 19556 14876 19612
rect 14812 19552 14876 19556
rect 14892 19612 14956 19616
rect 14892 19556 14896 19612
rect 14896 19556 14952 19612
rect 14952 19556 14956 19612
rect 14892 19552 14956 19556
rect 14972 19612 15036 19616
rect 14972 19556 14976 19612
rect 14976 19556 15032 19612
rect 15032 19556 15036 19612
rect 14972 19552 15036 19556
rect 20652 19612 20716 19616
rect 20652 19556 20656 19612
rect 20656 19556 20712 19612
rect 20712 19556 20716 19612
rect 20652 19552 20716 19556
rect 20732 19612 20796 19616
rect 20732 19556 20736 19612
rect 20736 19556 20792 19612
rect 20792 19556 20796 19612
rect 20732 19552 20796 19556
rect 20812 19612 20876 19616
rect 20812 19556 20816 19612
rect 20816 19556 20872 19612
rect 20872 19556 20876 19612
rect 20812 19552 20876 19556
rect 20892 19612 20956 19616
rect 20892 19556 20896 19612
rect 20896 19556 20952 19612
rect 20952 19556 20956 19612
rect 20892 19552 20956 19556
rect 20972 19612 21036 19616
rect 20972 19556 20976 19612
rect 20976 19556 21032 19612
rect 21032 19556 21036 19612
rect 20972 19552 21036 19556
rect 1912 19068 1976 19072
rect 1912 19012 1916 19068
rect 1916 19012 1972 19068
rect 1972 19012 1976 19068
rect 1912 19008 1976 19012
rect 1992 19068 2056 19072
rect 1992 19012 1996 19068
rect 1996 19012 2052 19068
rect 2052 19012 2056 19068
rect 1992 19008 2056 19012
rect 2072 19068 2136 19072
rect 2072 19012 2076 19068
rect 2076 19012 2132 19068
rect 2132 19012 2136 19068
rect 2072 19008 2136 19012
rect 2152 19068 2216 19072
rect 2152 19012 2156 19068
rect 2156 19012 2212 19068
rect 2212 19012 2216 19068
rect 2152 19008 2216 19012
rect 2232 19068 2296 19072
rect 2232 19012 2236 19068
rect 2236 19012 2292 19068
rect 2292 19012 2296 19068
rect 2232 19008 2296 19012
rect 7912 19068 7976 19072
rect 7912 19012 7916 19068
rect 7916 19012 7972 19068
rect 7972 19012 7976 19068
rect 7912 19008 7976 19012
rect 7992 19068 8056 19072
rect 7992 19012 7996 19068
rect 7996 19012 8052 19068
rect 8052 19012 8056 19068
rect 7992 19008 8056 19012
rect 8072 19068 8136 19072
rect 8072 19012 8076 19068
rect 8076 19012 8132 19068
rect 8132 19012 8136 19068
rect 8072 19008 8136 19012
rect 8152 19068 8216 19072
rect 8152 19012 8156 19068
rect 8156 19012 8212 19068
rect 8212 19012 8216 19068
rect 8152 19008 8216 19012
rect 8232 19068 8296 19072
rect 8232 19012 8236 19068
rect 8236 19012 8292 19068
rect 8292 19012 8296 19068
rect 8232 19008 8296 19012
rect 13912 19068 13976 19072
rect 13912 19012 13916 19068
rect 13916 19012 13972 19068
rect 13972 19012 13976 19068
rect 13912 19008 13976 19012
rect 13992 19068 14056 19072
rect 13992 19012 13996 19068
rect 13996 19012 14052 19068
rect 14052 19012 14056 19068
rect 13992 19008 14056 19012
rect 14072 19068 14136 19072
rect 14072 19012 14076 19068
rect 14076 19012 14132 19068
rect 14132 19012 14136 19068
rect 14072 19008 14136 19012
rect 14152 19068 14216 19072
rect 14152 19012 14156 19068
rect 14156 19012 14212 19068
rect 14212 19012 14216 19068
rect 14152 19008 14216 19012
rect 14232 19068 14296 19072
rect 14232 19012 14236 19068
rect 14236 19012 14292 19068
rect 14292 19012 14296 19068
rect 14232 19008 14296 19012
rect 19912 19068 19976 19072
rect 19912 19012 19916 19068
rect 19916 19012 19972 19068
rect 19972 19012 19976 19068
rect 19912 19008 19976 19012
rect 19992 19068 20056 19072
rect 19992 19012 19996 19068
rect 19996 19012 20052 19068
rect 20052 19012 20056 19068
rect 19992 19008 20056 19012
rect 20072 19068 20136 19072
rect 20072 19012 20076 19068
rect 20076 19012 20132 19068
rect 20132 19012 20136 19068
rect 20072 19008 20136 19012
rect 20152 19068 20216 19072
rect 20152 19012 20156 19068
rect 20156 19012 20212 19068
rect 20212 19012 20216 19068
rect 20152 19008 20216 19012
rect 20232 19068 20296 19072
rect 20232 19012 20236 19068
rect 20236 19012 20292 19068
rect 20292 19012 20296 19068
rect 20232 19008 20296 19012
rect 2652 18524 2716 18528
rect 2652 18468 2656 18524
rect 2656 18468 2712 18524
rect 2712 18468 2716 18524
rect 2652 18464 2716 18468
rect 2732 18524 2796 18528
rect 2732 18468 2736 18524
rect 2736 18468 2792 18524
rect 2792 18468 2796 18524
rect 2732 18464 2796 18468
rect 2812 18524 2876 18528
rect 2812 18468 2816 18524
rect 2816 18468 2872 18524
rect 2872 18468 2876 18524
rect 2812 18464 2876 18468
rect 2892 18524 2956 18528
rect 2892 18468 2896 18524
rect 2896 18468 2952 18524
rect 2952 18468 2956 18524
rect 2892 18464 2956 18468
rect 2972 18524 3036 18528
rect 2972 18468 2976 18524
rect 2976 18468 3032 18524
rect 3032 18468 3036 18524
rect 2972 18464 3036 18468
rect 8652 18524 8716 18528
rect 8652 18468 8656 18524
rect 8656 18468 8712 18524
rect 8712 18468 8716 18524
rect 8652 18464 8716 18468
rect 8732 18524 8796 18528
rect 8732 18468 8736 18524
rect 8736 18468 8792 18524
rect 8792 18468 8796 18524
rect 8732 18464 8796 18468
rect 8812 18524 8876 18528
rect 8812 18468 8816 18524
rect 8816 18468 8872 18524
rect 8872 18468 8876 18524
rect 8812 18464 8876 18468
rect 8892 18524 8956 18528
rect 8892 18468 8896 18524
rect 8896 18468 8952 18524
rect 8952 18468 8956 18524
rect 8892 18464 8956 18468
rect 8972 18524 9036 18528
rect 8972 18468 8976 18524
rect 8976 18468 9032 18524
rect 9032 18468 9036 18524
rect 8972 18464 9036 18468
rect 14652 18524 14716 18528
rect 14652 18468 14656 18524
rect 14656 18468 14712 18524
rect 14712 18468 14716 18524
rect 14652 18464 14716 18468
rect 14732 18524 14796 18528
rect 14732 18468 14736 18524
rect 14736 18468 14792 18524
rect 14792 18468 14796 18524
rect 14732 18464 14796 18468
rect 14812 18524 14876 18528
rect 14812 18468 14816 18524
rect 14816 18468 14872 18524
rect 14872 18468 14876 18524
rect 14812 18464 14876 18468
rect 14892 18524 14956 18528
rect 14892 18468 14896 18524
rect 14896 18468 14952 18524
rect 14952 18468 14956 18524
rect 14892 18464 14956 18468
rect 14972 18524 15036 18528
rect 14972 18468 14976 18524
rect 14976 18468 15032 18524
rect 15032 18468 15036 18524
rect 14972 18464 15036 18468
rect 20652 18524 20716 18528
rect 20652 18468 20656 18524
rect 20656 18468 20712 18524
rect 20712 18468 20716 18524
rect 20652 18464 20716 18468
rect 20732 18524 20796 18528
rect 20732 18468 20736 18524
rect 20736 18468 20792 18524
rect 20792 18468 20796 18524
rect 20732 18464 20796 18468
rect 20812 18524 20876 18528
rect 20812 18468 20816 18524
rect 20816 18468 20872 18524
rect 20872 18468 20876 18524
rect 20812 18464 20876 18468
rect 20892 18524 20956 18528
rect 20892 18468 20896 18524
rect 20896 18468 20952 18524
rect 20952 18468 20956 18524
rect 20892 18464 20956 18468
rect 20972 18524 21036 18528
rect 20972 18468 20976 18524
rect 20976 18468 21032 18524
rect 21032 18468 21036 18524
rect 20972 18464 21036 18468
rect 1912 17980 1976 17984
rect 1912 17924 1916 17980
rect 1916 17924 1972 17980
rect 1972 17924 1976 17980
rect 1912 17920 1976 17924
rect 1992 17980 2056 17984
rect 1992 17924 1996 17980
rect 1996 17924 2052 17980
rect 2052 17924 2056 17980
rect 1992 17920 2056 17924
rect 2072 17980 2136 17984
rect 2072 17924 2076 17980
rect 2076 17924 2132 17980
rect 2132 17924 2136 17980
rect 2072 17920 2136 17924
rect 2152 17980 2216 17984
rect 2152 17924 2156 17980
rect 2156 17924 2212 17980
rect 2212 17924 2216 17980
rect 2152 17920 2216 17924
rect 2232 17980 2296 17984
rect 2232 17924 2236 17980
rect 2236 17924 2292 17980
rect 2292 17924 2296 17980
rect 2232 17920 2296 17924
rect 7912 17980 7976 17984
rect 7912 17924 7916 17980
rect 7916 17924 7972 17980
rect 7972 17924 7976 17980
rect 7912 17920 7976 17924
rect 7992 17980 8056 17984
rect 7992 17924 7996 17980
rect 7996 17924 8052 17980
rect 8052 17924 8056 17980
rect 7992 17920 8056 17924
rect 8072 17980 8136 17984
rect 8072 17924 8076 17980
rect 8076 17924 8132 17980
rect 8132 17924 8136 17980
rect 8072 17920 8136 17924
rect 8152 17980 8216 17984
rect 8152 17924 8156 17980
rect 8156 17924 8212 17980
rect 8212 17924 8216 17980
rect 8152 17920 8216 17924
rect 8232 17980 8296 17984
rect 8232 17924 8236 17980
rect 8236 17924 8292 17980
rect 8292 17924 8296 17980
rect 8232 17920 8296 17924
rect 13912 17980 13976 17984
rect 13912 17924 13916 17980
rect 13916 17924 13972 17980
rect 13972 17924 13976 17980
rect 13912 17920 13976 17924
rect 13992 17980 14056 17984
rect 13992 17924 13996 17980
rect 13996 17924 14052 17980
rect 14052 17924 14056 17980
rect 13992 17920 14056 17924
rect 14072 17980 14136 17984
rect 14072 17924 14076 17980
rect 14076 17924 14132 17980
rect 14132 17924 14136 17980
rect 14072 17920 14136 17924
rect 14152 17980 14216 17984
rect 14152 17924 14156 17980
rect 14156 17924 14212 17980
rect 14212 17924 14216 17980
rect 14152 17920 14216 17924
rect 14232 17980 14296 17984
rect 14232 17924 14236 17980
rect 14236 17924 14292 17980
rect 14292 17924 14296 17980
rect 14232 17920 14296 17924
rect 19912 17980 19976 17984
rect 19912 17924 19916 17980
rect 19916 17924 19972 17980
rect 19972 17924 19976 17980
rect 19912 17920 19976 17924
rect 19992 17980 20056 17984
rect 19992 17924 19996 17980
rect 19996 17924 20052 17980
rect 20052 17924 20056 17980
rect 19992 17920 20056 17924
rect 20072 17980 20136 17984
rect 20072 17924 20076 17980
rect 20076 17924 20132 17980
rect 20132 17924 20136 17980
rect 20072 17920 20136 17924
rect 20152 17980 20216 17984
rect 20152 17924 20156 17980
rect 20156 17924 20212 17980
rect 20212 17924 20216 17980
rect 20152 17920 20216 17924
rect 20232 17980 20296 17984
rect 20232 17924 20236 17980
rect 20236 17924 20292 17980
rect 20292 17924 20296 17980
rect 20232 17920 20296 17924
rect 2652 17436 2716 17440
rect 2652 17380 2656 17436
rect 2656 17380 2712 17436
rect 2712 17380 2716 17436
rect 2652 17376 2716 17380
rect 2732 17436 2796 17440
rect 2732 17380 2736 17436
rect 2736 17380 2792 17436
rect 2792 17380 2796 17436
rect 2732 17376 2796 17380
rect 2812 17436 2876 17440
rect 2812 17380 2816 17436
rect 2816 17380 2872 17436
rect 2872 17380 2876 17436
rect 2812 17376 2876 17380
rect 2892 17436 2956 17440
rect 2892 17380 2896 17436
rect 2896 17380 2952 17436
rect 2952 17380 2956 17436
rect 2892 17376 2956 17380
rect 2972 17436 3036 17440
rect 2972 17380 2976 17436
rect 2976 17380 3032 17436
rect 3032 17380 3036 17436
rect 2972 17376 3036 17380
rect 8652 17436 8716 17440
rect 8652 17380 8656 17436
rect 8656 17380 8712 17436
rect 8712 17380 8716 17436
rect 8652 17376 8716 17380
rect 8732 17436 8796 17440
rect 8732 17380 8736 17436
rect 8736 17380 8792 17436
rect 8792 17380 8796 17436
rect 8732 17376 8796 17380
rect 8812 17436 8876 17440
rect 8812 17380 8816 17436
rect 8816 17380 8872 17436
rect 8872 17380 8876 17436
rect 8812 17376 8876 17380
rect 8892 17436 8956 17440
rect 8892 17380 8896 17436
rect 8896 17380 8952 17436
rect 8952 17380 8956 17436
rect 8892 17376 8956 17380
rect 8972 17436 9036 17440
rect 8972 17380 8976 17436
rect 8976 17380 9032 17436
rect 9032 17380 9036 17436
rect 8972 17376 9036 17380
rect 14652 17436 14716 17440
rect 14652 17380 14656 17436
rect 14656 17380 14712 17436
rect 14712 17380 14716 17436
rect 14652 17376 14716 17380
rect 14732 17436 14796 17440
rect 14732 17380 14736 17436
rect 14736 17380 14792 17436
rect 14792 17380 14796 17436
rect 14732 17376 14796 17380
rect 14812 17436 14876 17440
rect 14812 17380 14816 17436
rect 14816 17380 14872 17436
rect 14872 17380 14876 17436
rect 14812 17376 14876 17380
rect 14892 17436 14956 17440
rect 14892 17380 14896 17436
rect 14896 17380 14952 17436
rect 14952 17380 14956 17436
rect 14892 17376 14956 17380
rect 14972 17436 15036 17440
rect 14972 17380 14976 17436
rect 14976 17380 15032 17436
rect 15032 17380 15036 17436
rect 14972 17376 15036 17380
rect 20652 17436 20716 17440
rect 20652 17380 20656 17436
rect 20656 17380 20712 17436
rect 20712 17380 20716 17436
rect 20652 17376 20716 17380
rect 20732 17436 20796 17440
rect 20732 17380 20736 17436
rect 20736 17380 20792 17436
rect 20792 17380 20796 17436
rect 20732 17376 20796 17380
rect 20812 17436 20876 17440
rect 20812 17380 20816 17436
rect 20816 17380 20872 17436
rect 20872 17380 20876 17436
rect 20812 17376 20876 17380
rect 20892 17436 20956 17440
rect 20892 17380 20896 17436
rect 20896 17380 20952 17436
rect 20952 17380 20956 17436
rect 20892 17376 20956 17380
rect 20972 17436 21036 17440
rect 20972 17380 20976 17436
rect 20976 17380 21032 17436
rect 21032 17380 21036 17436
rect 20972 17376 21036 17380
rect 1912 16892 1976 16896
rect 1912 16836 1916 16892
rect 1916 16836 1972 16892
rect 1972 16836 1976 16892
rect 1912 16832 1976 16836
rect 1992 16892 2056 16896
rect 1992 16836 1996 16892
rect 1996 16836 2052 16892
rect 2052 16836 2056 16892
rect 1992 16832 2056 16836
rect 2072 16892 2136 16896
rect 2072 16836 2076 16892
rect 2076 16836 2132 16892
rect 2132 16836 2136 16892
rect 2072 16832 2136 16836
rect 2152 16892 2216 16896
rect 2152 16836 2156 16892
rect 2156 16836 2212 16892
rect 2212 16836 2216 16892
rect 2152 16832 2216 16836
rect 2232 16892 2296 16896
rect 2232 16836 2236 16892
rect 2236 16836 2292 16892
rect 2292 16836 2296 16892
rect 2232 16832 2296 16836
rect 7912 16892 7976 16896
rect 7912 16836 7916 16892
rect 7916 16836 7972 16892
rect 7972 16836 7976 16892
rect 7912 16832 7976 16836
rect 7992 16892 8056 16896
rect 7992 16836 7996 16892
rect 7996 16836 8052 16892
rect 8052 16836 8056 16892
rect 7992 16832 8056 16836
rect 8072 16892 8136 16896
rect 8072 16836 8076 16892
rect 8076 16836 8132 16892
rect 8132 16836 8136 16892
rect 8072 16832 8136 16836
rect 8152 16892 8216 16896
rect 8152 16836 8156 16892
rect 8156 16836 8212 16892
rect 8212 16836 8216 16892
rect 8152 16832 8216 16836
rect 8232 16892 8296 16896
rect 8232 16836 8236 16892
rect 8236 16836 8292 16892
rect 8292 16836 8296 16892
rect 8232 16832 8296 16836
rect 13912 16892 13976 16896
rect 13912 16836 13916 16892
rect 13916 16836 13972 16892
rect 13972 16836 13976 16892
rect 13912 16832 13976 16836
rect 13992 16892 14056 16896
rect 13992 16836 13996 16892
rect 13996 16836 14052 16892
rect 14052 16836 14056 16892
rect 13992 16832 14056 16836
rect 14072 16892 14136 16896
rect 14072 16836 14076 16892
rect 14076 16836 14132 16892
rect 14132 16836 14136 16892
rect 14072 16832 14136 16836
rect 14152 16892 14216 16896
rect 14152 16836 14156 16892
rect 14156 16836 14212 16892
rect 14212 16836 14216 16892
rect 14152 16832 14216 16836
rect 14232 16892 14296 16896
rect 14232 16836 14236 16892
rect 14236 16836 14292 16892
rect 14292 16836 14296 16892
rect 14232 16832 14296 16836
rect 19912 16892 19976 16896
rect 19912 16836 19916 16892
rect 19916 16836 19972 16892
rect 19972 16836 19976 16892
rect 19912 16832 19976 16836
rect 19992 16892 20056 16896
rect 19992 16836 19996 16892
rect 19996 16836 20052 16892
rect 20052 16836 20056 16892
rect 19992 16832 20056 16836
rect 20072 16892 20136 16896
rect 20072 16836 20076 16892
rect 20076 16836 20132 16892
rect 20132 16836 20136 16892
rect 20072 16832 20136 16836
rect 20152 16892 20216 16896
rect 20152 16836 20156 16892
rect 20156 16836 20212 16892
rect 20212 16836 20216 16892
rect 20152 16832 20216 16836
rect 20232 16892 20296 16896
rect 20232 16836 20236 16892
rect 20236 16836 20292 16892
rect 20292 16836 20296 16892
rect 20232 16832 20296 16836
rect 2652 16348 2716 16352
rect 2652 16292 2656 16348
rect 2656 16292 2712 16348
rect 2712 16292 2716 16348
rect 2652 16288 2716 16292
rect 2732 16348 2796 16352
rect 2732 16292 2736 16348
rect 2736 16292 2792 16348
rect 2792 16292 2796 16348
rect 2732 16288 2796 16292
rect 2812 16348 2876 16352
rect 2812 16292 2816 16348
rect 2816 16292 2872 16348
rect 2872 16292 2876 16348
rect 2812 16288 2876 16292
rect 2892 16348 2956 16352
rect 2892 16292 2896 16348
rect 2896 16292 2952 16348
rect 2952 16292 2956 16348
rect 2892 16288 2956 16292
rect 2972 16348 3036 16352
rect 2972 16292 2976 16348
rect 2976 16292 3032 16348
rect 3032 16292 3036 16348
rect 2972 16288 3036 16292
rect 8652 16348 8716 16352
rect 8652 16292 8656 16348
rect 8656 16292 8712 16348
rect 8712 16292 8716 16348
rect 8652 16288 8716 16292
rect 8732 16348 8796 16352
rect 8732 16292 8736 16348
rect 8736 16292 8792 16348
rect 8792 16292 8796 16348
rect 8732 16288 8796 16292
rect 8812 16348 8876 16352
rect 8812 16292 8816 16348
rect 8816 16292 8872 16348
rect 8872 16292 8876 16348
rect 8812 16288 8876 16292
rect 8892 16348 8956 16352
rect 8892 16292 8896 16348
rect 8896 16292 8952 16348
rect 8952 16292 8956 16348
rect 8892 16288 8956 16292
rect 8972 16348 9036 16352
rect 8972 16292 8976 16348
rect 8976 16292 9032 16348
rect 9032 16292 9036 16348
rect 8972 16288 9036 16292
rect 14652 16348 14716 16352
rect 14652 16292 14656 16348
rect 14656 16292 14712 16348
rect 14712 16292 14716 16348
rect 14652 16288 14716 16292
rect 14732 16348 14796 16352
rect 14732 16292 14736 16348
rect 14736 16292 14792 16348
rect 14792 16292 14796 16348
rect 14732 16288 14796 16292
rect 14812 16348 14876 16352
rect 14812 16292 14816 16348
rect 14816 16292 14872 16348
rect 14872 16292 14876 16348
rect 14812 16288 14876 16292
rect 14892 16348 14956 16352
rect 14892 16292 14896 16348
rect 14896 16292 14952 16348
rect 14952 16292 14956 16348
rect 14892 16288 14956 16292
rect 14972 16348 15036 16352
rect 14972 16292 14976 16348
rect 14976 16292 15032 16348
rect 15032 16292 15036 16348
rect 14972 16288 15036 16292
rect 20652 16348 20716 16352
rect 20652 16292 20656 16348
rect 20656 16292 20712 16348
rect 20712 16292 20716 16348
rect 20652 16288 20716 16292
rect 20732 16348 20796 16352
rect 20732 16292 20736 16348
rect 20736 16292 20792 16348
rect 20792 16292 20796 16348
rect 20732 16288 20796 16292
rect 20812 16348 20876 16352
rect 20812 16292 20816 16348
rect 20816 16292 20872 16348
rect 20872 16292 20876 16348
rect 20812 16288 20876 16292
rect 20892 16348 20956 16352
rect 20892 16292 20896 16348
rect 20896 16292 20952 16348
rect 20952 16292 20956 16348
rect 20892 16288 20956 16292
rect 20972 16348 21036 16352
rect 20972 16292 20976 16348
rect 20976 16292 21032 16348
rect 21032 16292 21036 16348
rect 20972 16288 21036 16292
rect 1912 15804 1976 15808
rect 1912 15748 1916 15804
rect 1916 15748 1972 15804
rect 1972 15748 1976 15804
rect 1912 15744 1976 15748
rect 1992 15804 2056 15808
rect 1992 15748 1996 15804
rect 1996 15748 2052 15804
rect 2052 15748 2056 15804
rect 1992 15744 2056 15748
rect 2072 15804 2136 15808
rect 2072 15748 2076 15804
rect 2076 15748 2132 15804
rect 2132 15748 2136 15804
rect 2072 15744 2136 15748
rect 2152 15804 2216 15808
rect 2152 15748 2156 15804
rect 2156 15748 2212 15804
rect 2212 15748 2216 15804
rect 2152 15744 2216 15748
rect 2232 15804 2296 15808
rect 2232 15748 2236 15804
rect 2236 15748 2292 15804
rect 2292 15748 2296 15804
rect 2232 15744 2296 15748
rect 7912 15804 7976 15808
rect 7912 15748 7916 15804
rect 7916 15748 7972 15804
rect 7972 15748 7976 15804
rect 7912 15744 7976 15748
rect 7992 15804 8056 15808
rect 7992 15748 7996 15804
rect 7996 15748 8052 15804
rect 8052 15748 8056 15804
rect 7992 15744 8056 15748
rect 8072 15804 8136 15808
rect 8072 15748 8076 15804
rect 8076 15748 8132 15804
rect 8132 15748 8136 15804
rect 8072 15744 8136 15748
rect 8152 15804 8216 15808
rect 8152 15748 8156 15804
rect 8156 15748 8212 15804
rect 8212 15748 8216 15804
rect 8152 15744 8216 15748
rect 8232 15804 8296 15808
rect 8232 15748 8236 15804
rect 8236 15748 8292 15804
rect 8292 15748 8296 15804
rect 8232 15744 8296 15748
rect 13912 15804 13976 15808
rect 13912 15748 13916 15804
rect 13916 15748 13972 15804
rect 13972 15748 13976 15804
rect 13912 15744 13976 15748
rect 13992 15804 14056 15808
rect 13992 15748 13996 15804
rect 13996 15748 14052 15804
rect 14052 15748 14056 15804
rect 13992 15744 14056 15748
rect 14072 15804 14136 15808
rect 14072 15748 14076 15804
rect 14076 15748 14132 15804
rect 14132 15748 14136 15804
rect 14072 15744 14136 15748
rect 14152 15804 14216 15808
rect 14152 15748 14156 15804
rect 14156 15748 14212 15804
rect 14212 15748 14216 15804
rect 14152 15744 14216 15748
rect 14232 15804 14296 15808
rect 14232 15748 14236 15804
rect 14236 15748 14292 15804
rect 14292 15748 14296 15804
rect 14232 15744 14296 15748
rect 19912 15804 19976 15808
rect 19912 15748 19916 15804
rect 19916 15748 19972 15804
rect 19972 15748 19976 15804
rect 19912 15744 19976 15748
rect 19992 15804 20056 15808
rect 19992 15748 19996 15804
rect 19996 15748 20052 15804
rect 20052 15748 20056 15804
rect 19992 15744 20056 15748
rect 20072 15804 20136 15808
rect 20072 15748 20076 15804
rect 20076 15748 20132 15804
rect 20132 15748 20136 15804
rect 20072 15744 20136 15748
rect 20152 15804 20216 15808
rect 20152 15748 20156 15804
rect 20156 15748 20212 15804
rect 20212 15748 20216 15804
rect 20152 15744 20216 15748
rect 20232 15804 20296 15808
rect 20232 15748 20236 15804
rect 20236 15748 20292 15804
rect 20292 15748 20296 15804
rect 20232 15744 20296 15748
rect 2652 15260 2716 15264
rect 2652 15204 2656 15260
rect 2656 15204 2712 15260
rect 2712 15204 2716 15260
rect 2652 15200 2716 15204
rect 2732 15260 2796 15264
rect 2732 15204 2736 15260
rect 2736 15204 2792 15260
rect 2792 15204 2796 15260
rect 2732 15200 2796 15204
rect 2812 15260 2876 15264
rect 2812 15204 2816 15260
rect 2816 15204 2872 15260
rect 2872 15204 2876 15260
rect 2812 15200 2876 15204
rect 2892 15260 2956 15264
rect 2892 15204 2896 15260
rect 2896 15204 2952 15260
rect 2952 15204 2956 15260
rect 2892 15200 2956 15204
rect 2972 15260 3036 15264
rect 2972 15204 2976 15260
rect 2976 15204 3032 15260
rect 3032 15204 3036 15260
rect 2972 15200 3036 15204
rect 8652 15260 8716 15264
rect 8652 15204 8656 15260
rect 8656 15204 8712 15260
rect 8712 15204 8716 15260
rect 8652 15200 8716 15204
rect 8732 15260 8796 15264
rect 8732 15204 8736 15260
rect 8736 15204 8792 15260
rect 8792 15204 8796 15260
rect 8732 15200 8796 15204
rect 8812 15260 8876 15264
rect 8812 15204 8816 15260
rect 8816 15204 8872 15260
rect 8872 15204 8876 15260
rect 8812 15200 8876 15204
rect 8892 15260 8956 15264
rect 8892 15204 8896 15260
rect 8896 15204 8952 15260
rect 8952 15204 8956 15260
rect 8892 15200 8956 15204
rect 8972 15260 9036 15264
rect 8972 15204 8976 15260
rect 8976 15204 9032 15260
rect 9032 15204 9036 15260
rect 8972 15200 9036 15204
rect 14652 15260 14716 15264
rect 14652 15204 14656 15260
rect 14656 15204 14712 15260
rect 14712 15204 14716 15260
rect 14652 15200 14716 15204
rect 14732 15260 14796 15264
rect 14732 15204 14736 15260
rect 14736 15204 14792 15260
rect 14792 15204 14796 15260
rect 14732 15200 14796 15204
rect 14812 15260 14876 15264
rect 14812 15204 14816 15260
rect 14816 15204 14872 15260
rect 14872 15204 14876 15260
rect 14812 15200 14876 15204
rect 14892 15260 14956 15264
rect 14892 15204 14896 15260
rect 14896 15204 14952 15260
rect 14952 15204 14956 15260
rect 14892 15200 14956 15204
rect 14972 15260 15036 15264
rect 14972 15204 14976 15260
rect 14976 15204 15032 15260
rect 15032 15204 15036 15260
rect 14972 15200 15036 15204
rect 20652 15260 20716 15264
rect 20652 15204 20656 15260
rect 20656 15204 20712 15260
rect 20712 15204 20716 15260
rect 20652 15200 20716 15204
rect 20732 15260 20796 15264
rect 20732 15204 20736 15260
rect 20736 15204 20792 15260
rect 20792 15204 20796 15260
rect 20732 15200 20796 15204
rect 20812 15260 20876 15264
rect 20812 15204 20816 15260
rect 20816 15204 20872 15260
rect 20872 15204 20876 15260
rect 20812 15200 20876 15204
rect 20892 15260 20956 15264
rect 20892 15204 20896 15260
rect 20896 15204 20952 15260
rect 20952 15204 20956 15260
rect 20892 15200 20956 15204
rect 20972 15260 21036 15264
rect 20972 15204 20976 15260
rect 20976 15204 21032 15260
rect 21032 15204 21036 15260
rect 20972 15200 21036 15204
rect 1912 14716 1976 14720
rect 1912 14660 1916 14716
rect 1916 14660 1972 14716
rect 1972 14660 1976 14716
rect 1912 14656 1976 14660
rect 1992 14716 2056 14720
rect 1992 14660 1996 14716
rect 1996 14660 2052 14716
rect 2052 14660 2056 14716
rect 1992 14656 2056 14660
rect 2072 14716 2136 14720
rect 2072 14660 2076 14716
rect 2076 14660 2132 14716
rect 2132 14660 2136 14716
rect 2072 14656 2136 14660
rect 2152 14716 2216 14720
rect 2152 14660 2156 14716
rect 2156 14660 2212 14716
rect 2212 14660 2216 14716
rect 2152 14656 2216 14660
rect 2232 14716 2296 14720
rect 2232 14660 2236 14716
rect 2236 14660 2292 14716
rect 2292 14660 2296 14716
rect 2232 14656 2296 14660
rect 7912 14716 7976 14720
rect 7912 14660 7916 14716
rect 7916 14660 7972 14716
rect 7972 14660 7976 14716
rect 7912 14656 7976 14660
rect 7992 14716 8056 14720
rect 7992 14660 7996 14716
rect 7996 14660 8052 14716
rect 8052 14660 8056 14716
rect 7992 14656 8056 14660
rect 8072 14716 8136 14720
rect 8072 14660 8076 14716
rect 8076 14660 8132 14716
rect 8132 14660 8136 14716
rect 8072 14656 8136 14660
rect 8152 14716 8216 14720
rect 8152 14660 8156 14716
rect 8156 14660 8212 14716
rect 8212 14660 8216 14716
rect 8152 14656 8216 14660
rect 8232 14716 8296 14720
rect 8232 14660 8236 14716
rect 8236 14660 8292 14716
rect 8292 14660 8296 14716
rect 8232 14656 8296 14660
rect 13912 14716 13976 14720
rect 13912 14660 13916 14716
rect 13916 14660 13972 14716
rect 13972 14660 13976 14716
rect 13912 14656 13976 14660
rect 13992 14716 14056 14720
rect 13992 14660 13996 14716
rect 13996 14660 14052 14716
rect 14052 14660 14056 14716
rect 13992 14656 14056 14660
rect 14072 14716 14136 14720
rect 14072 14660 14076 14716
rect 14076 14660 14132 14716
rect 14132 14660 14136 14716
rect 14072 14656 14136 14660
rect 14152 14716 14216 14720
rect 14152 14660 14156 14716
rect 14156 14660 14212 14716
rect 14212 14660 14216 14716
rect 14152 14656 14216 14660
rect 14232 14716 14296 14720
rect 14232 14660 14236 14716
rect 14236 14660 14292 14716
rect 14292 14660 14296 14716
rect 14232 14656 14296 14660
rect 19912 14716 19976 14720
rect 19912 14660 19916 14716
rect 19916 14660 19972 14716
rect 19972 14660 19976 14716
rect 19912 14656 19976 14660
rect 19992 14716 20056 14720
rect 19992 14660 19996 14716
rect 19996 14660 20052 14716
rect 20052 14660 20056 14716
rect 19992 14656 20056 14660
rect 20072 14716 20136 14720
rect 20072 14660 20076 14716
rect 20076 14660 20132 14716
rect 20132 14660 20136 14716
rect 20072 14656 20136 14660
rect 20152 14716 20216 14720
rect 20152 14660 20156 14716
rect 20156 14660 20212 14716
rect 20212 14660 20216 14716
rect 20152 14656 20216 14660
rect 20232 14716 20296 14720
rect 20232 14660 20236 14716
rect 20236 14660 20292 14716
rect 20292 14660 20296 14716
rect 20232 14656 20296 14660
rect 2652 14172 2716 14176
rect 2652 14116 2656 14172
rect 2656 14116 2712 14172
rect 2712 14116 2716 14172
rect 2652 14112 2716 14116
rect 2732 14172 2796 14176
rect 2732 14116 2736 14172
rect 2736 14116 2792 14172
rect 2792 14116 2796 14172
rect 2732 14112 2796 14116
rect 2812 14172 2876 14176
rect 2812 14116 2816 14172
rect 2816 14116 2872 14172
rect 2872 14116 2876 14172
rect 2812 14112 2876 14116
rect 2892 14172 2956 14176
rect 2892 14116 2896 14172
rect 2896 14116 2952 14172
rect 2952 14116 2956 14172
rect 2892 14112 2956 14116
rect 2972 14172 3036 14176
rect 2972 14116 2976 14172
rect 2976 14116 3032 14172
rect 3032 14116 3036 14172
rect 2972 14112 3036 14116
rect 8652 14172 8716 14176
rect 8652 14116 8656 14172
rect 8656 14116 8712 14172
rect 8712 14116 8716 14172
rect 8652 14112 8716 14116
rect 8732 14172 8796 14176
rect 8732 14116 8736 14172
rect 8736 14116 8792 14172
rect 8792 14116 8796 14172
rect 8732 14112 8796 14116
rect 8812 14172 8876 14176
rect 8812 14116 8816 14172
rect 8816 14116 8872 14172
rect 8872 14116 8876 14172
rect 8812 14112 8876 14116
rect 8892 14172 8956 14176
rect 8892 14116 8896 14172
rect 8896 14116 8952 14172
rect 8952 14116 8956 14172
rect 8892 14112 8956 14116
rect 8972 14172 9036 14176
rect 8972 14116 8976 14172
rect 8976 14116 9032 14172
rect 9032 14116 9036 14172
rect 8972 14112 9036 14116
rect 14652 14172 14716 14176
rect 14652 14116 14656 14172
rect 14656 14116 14712 14172
rect 14712 14116 14716 14172
rect 14652 14112 14716 14116
rect 14732 14172 14796 14176
rect 14732 14116 14736 14172
rect 14736 14116 14792 14172
rect 14792 14116 14796 14172
rect 14732 14112 14796 14116
rect 14812 14172 14876 14176
rect 14812 14116 14816 14172
rect 14816 14116 14872 14172
rect 14872 14116 14876 14172
rect 14812 14112 14876 14116
rect 14892 14172 14956 14176
rect 14892 14116 14896 14172
rect 14896 14116 14952 14172
rect 14952 14116 14956 14172
rect 14892 14112 14956 14116
rect 14972 14172 15036 14176
rect 14972 14116 14976 14172
rect 14976 14116 15032 14172
rect 15032 14116 15036 14172
rect 14972 14112 15036 14116
rect 20652 14172 20716 14176
rect 20652 14116 20656 14172
rect 20656 14116 20712 14172
rect 20712 14116 20716 14172
rect 20652 14112 20716 14116
rect 20732 14172 20796 14176
rect 20732 14116 20736 14172
rect 20736 14116 20792 14172
rect 20792 14116 20796 14172
rect 20732 14112 20796 14116
rect 20812 14172 20876 14176
rect 20812 14116 20816 14172
rect 20816 14116 20872 14172
rect 20872 14116 20876 14172
rect 20812 14112 20876 14116
rect 20892 14172 20956 14176
rect 20892 14116 20896 14172
rect 20896 14116 20952 14172
rect 20952 14116 20956 14172
rect 20892 14112 20956 14116
rect 20972 14172 21036 14176
rect 20972 14116 20976 14172
rect 20976 14116 21032 14172
rect 21032 14116 21036 14172
rect 20972 14112 21036 14116
rect 1912 13628 1976 13632
rect 1912 13572 1916 13628
rect 1916 13572 1972 13628
rect 1972 13572 1976 13628
rect 1912 13568 1976 13572
rect 1992 13628 2056 13632
rect 1992 13572 1996 13628
rect 1996 13572 2052 13628
rect 2052 13572 2056 13628
rect 1992 13568 2056 13572
rect 2072 13628 2136 13632
rect 2072 13572 2076 13628
rect 2076 13572 2132 13628
rect 2132 13572 2136 13628
rect 2072 13568 2136 13572
rect 2152 13628 2216 13632
rect 2152 13572 2156 13628
rect 2156 13572 2212 13628
rect 2212 13572 2216 13628
rect 2152 13568 2216 13572
rect 2232 13628 2296 13632
rect 2232 13572 2236 13628
rect 2236 13572 2292 13628
rect 2292 13572 2296 13628
rect 2232 13568 2296 13572
rect 7912 13628 7976 13632
rect 7912 13572 7916 13628
rect 7916 13572 7972 13628
rect 7972 13572 7976 13628
rect 7912 13568 7976 13572
rect 7992 13628 8056 13632
rect 7992 13572 7996 13628
rect 7996 13572 8052 13628
rect 8052 13572 8056 13628
rect 7992 13568 8056 13572
rect 8072 13628 8136 13632
rect 8072 13572 8076 13628
rect 8076 13572 8132 13628
rect 8132 13572 8136 13628
rect 8072 13568 8136 13572
rect 8152 13628 8216 13632
rect 8152 13572 8156 13628
rect 8156 13572 8212 13628
rect 8212 13572 8216 13628
rect 8152 13568 8216 13572
rect 8232 13628 8296 13632
rect 8232 13572 8236 13628
rect 8236 13572 8292 13628
rect 8292 13572 8296 13628
rect 8232 13568 8296 13572
rect 13912 13628 13976 13632
rect 13912 13572 13916 13628
rect 13916 13572 13972 13628
rect 13972 13572 13976 13628
rect 13912 13568 13976 13572
rect 13992 13628 14056 13632
rect 13992 13572 13996 13628
rect 13996 13572 14052 13628
rect 14052 13572 14056 13628
rect 13992 13568 14056 13572
rect 14072 13628 14136 13632
rect 14072 13572 14076 13628
rect 14076 13572 14132 13628
rect 14132 13572 14136 13628
rect 14072 13568 14136 13572
rect 14152 13628 14216 13632
rect 14152 13572 14156 13628
rect 14156 13572 14212 13628
rect 14212 13572 14216 13628
rect 14152 13568 14216 13572
rect 14232 13628 14296 13632
rect 14232 13572 14236 13628
rect 14236 13572 14292 13628
rect 14292 13572 14296 13628
rect 14232 13568 14296 13572
rect 19912 13628 19976 13632
rect 19912 13572 19916 13628
rect 19916 13572 19972 13628
rect 19972 13572 19976 13628
rect 19912 13568 19976 13572
rect 19992 13628 20056 13632
rect 19992 13572 19996 13628
rect 19996 13572 20052 13628
rect 20052 13572 20056 13628
rect 19992 13568 20056 13572
rect 20072 13628 20136 13632
rect 20072 13572 20076 13628
rect 20076 13572 20132 13628
rect 20132 13572 20136 13628
rect 20072 13568 20136 13572
rect 20152 13628 20216 13632
rect 20152 13572 20156 13628
rect 20156 13572 20212 13628
rect 20212 13572 20216 13628
rect 20152 13568 20216 13572
rect 20232 13628 20296 13632
rect 20232 13572 20236 13628
rect 20236 13572 20292 13628
rect 20292 13572 20296 13628
rect 20232 13568 20296 13572
rect 2652 13084 2716 13088
rect 2652 13028 2656 13084
rect 2656 13028 2712 13084
rect 2712 13028 2716 13084
rect 2652 13024 2716 13028
rect 2732 13084 2796 13088
rect 2732 13028 2736 13084
rect 2736 13028 2792 13084
rect 2792 13028 2796 13084
rect 2732 13024 2796 13028
rect 2812 13084 2876 13088
rect 2812 13028 2816 13084
rect 2816 13028 2872 13084
rect 2872 13028 2876 13084
rect 2812 13024 2876 13028
rect 2892 13084 2956 13088
rect 2892 13028 2896 13084
rect 2896 13028 2952 13084
rect 2952 13028 2956 13084
rect 2892 13024 2956 13028
rect 2972 13084 3036 13088
rect 2972 13028 2976 13084
rect 2976 13028 3032 13084
rect 3032 13028 3036 13084
rect 2972 13024 3036 13028
rect 8652 13084 8716 13088
rect 8652 13028 8656 13084
rect 8656 13028 8712 13084
rect 8712 13028 8716 13084
rect 8652 13024 8716 13028
rect 8732 13084 8796 13088
rect 8732 13028 8736 13084
rect 8736 13028 8792 13084
rect 8792 13028 8796 13084
rect 8732 13024 8796 13028
rect 8812 13084 8876 13088
rect 8812 13028 8816 13084
rect 8816 13028 8872 13084
rect 8872 13028 8876 13084
rect 8812 13024 8876 13028
rect 8892 13084 8956 13088
rect 8892 13028 8896 13084
rect 8896 13028 8952 13084
rect 8952 13028 8956 13084
rect 8892 13024 8956 13028
rect 8972 13084 9036 13088
rect 8972 13028 8976 13084
rect 8976 13028 9032 13084
rect 9032 13028 9036 13084
rect 8972 13024 9036 13028
rect 14652 13084 14716 13088
rect 14652 13028 14656 13084
rect 14656 13028 14712 13084
rect 14712 13028 14716 13084
rect 14652 13024 14716 13028
rect 14732 13084 14796 13088
rect 14732 13028 14736 13084
rect 14736 13028 14792 13084
rect 14792 13028 14796 13084
rect 14732 13024 14796 13028
rect 14812 13084 14876 13088
rect 14812 13028 14816 13084
rect 14816 13028 14872 13084
rect 14872 13028 14876 13084
rect 14812 13024 14876 13028
rect 14892 13084 14956 13088
rect 14892 13028 14896 13084
rect 14896 13028 14952 13084
rect 14952 13028 14956 13084
rect 14892 13024 14956 13028
rect 14972 13084 15036 13088
rect 14972 13028 14976 13084
rect 14976 13028 15032 13084
rect 15032 13028 15036 13084
rect 14972 13024 15036 13028
rect 20652 13084 20716 13088
rect 20652 13028 20656 13084
rect 20656 13028 20712 13084
rect 20712 13028 20716 13084
rect 20652 13024 20716 13028
rect 20732 13084 20796 13088
rect 20732 13028 20736 13084
rect 20736 13028 20792 13084
rect 20792 13028 20796 13084
rect 20732 13024 20796 13028
rect 20812 13084 20876 13088
rect 20812 13028 20816 13084
rect 20816 13028 20872 13084
rect 20872 13028 20876 13084
rect 20812 13024 20876 13028
rect 20892 13084 20956 13088
rect 20892 13028 20896 13084
rect 20896 13028 20952 13084
rect 20952 13028 20956 13084
rect 20892 13024 20956 13028
rect 20972 13084 21036 13088
rect 20972 13028 20976 13084
rect 20976 13028 21032 13084
rect 21032 13028 21036 13084
rect 20972 13024 21036 13028
rect 9444 12744 9508 12748
rect 9444 12688 9458 12744
rect 9458 12688 9508 12744
rect 9444 12684 9508 12688
rect 1912 12540 1976 12544
rect 1912 12484 1916 12540
rect 1916 12484 1972 12540
rect 1972 12484 1976 12540
rect 1912 12480 1976 12484
rect 1992 12540 2056 12544
rect 1992 12484 1996 12540
rect 1996 12484 2052 12540
rect 2052 12484 2056 12540
rect 1992 12480 2056 12484
rect 2072 12540 2136 12544
rect 2072 12484 2076 12540
rect 2076 12484 2132 12540
rect 2132 12484 2136 12540
rect 2072 12480 2136 12484
rect 2152 12540 2216 12544
rect 2152 12484 2156 12540
rect 2156 12484 2212 12540
rect 2212 12484 2216 12540
rect 2152 12480 2216 12484
rect 2232 12540 2296 12544
rect 2232 12484 2236 12540
rect 2236 12484 2292 12540
rect 2292 12484 2296 12540
rect 2232 12480 2296 12484
rect 7912 12540 7976 12544
rect 7912 12484 7916 12540
rect 7916 12484 7972 12540
rect 7972 12484 7976 12540
rect 7912 12480 7976 12484
rect 7992 12540 8056 12544
rect 7992 12484 7996 12540
rect 7996 12484 8052 12540
rect 8052 12484 8056 12540
rect 7992 12480 8056 12484
rect 8072 12540 8136 12544
rect 8072 12484 8076 12540
rect 8076 12484 8132 12540
rect 8132 12484 8136 12540
rect 8072 12480 8136 12484
rect 8152 12540 8216 12544
rect 8152 12484 8156 12540
rect 8156 12484 8212 12540
rect 8212 12484 8216 12540
rect 8152 12480 8216 12484
rect 8232 12540 8296 12544
rect 8232 12484 8236 12540
rect 8236 12484 8292 12540
rect 8292 12484 8296 12540
rect 8232 12480 8296 12484
rect 13912 12540 13976 12544
rect 13912 12484 13916 12540
rect 13916 12484 13972 12540
rect 13972 12484 13976 12540
rect 13912 12480 13976 12484
rect 13992 12540 14056 12544
rect 13992 12484 13996 12540
rect 13996 12484 14052 12540
rect 14052 12484 14056 12540
rect 13992 12480 14056 12484
rect 14072 12540 14136 12544
rect 14072 12484 14076 12540
rect 14076 12484 14132 12540
rect 14132 12484 14136 12540
rect 14072 12480 14136 12484
rect 14152 12540 14216 12544
rect 14152 12484 14156 12540
rect 14156 12484 14212 12540
rect 14212 12484 14216 12540
rect 14152 12480 14216 12484
rect 14232 12540 14296 12544
rect 14232 12484 14236 12540
rect 14236 12484 14292 12540
rect 14292 12484 14296 12540
rect 14232 12480 14296 12484
rect 19912 12540 19976 12544
rect 19912 12484 19916 12540
rect 19916 12484 19972 12540
rect 19972 12484 19976 12540
rect 19912 12480 19976 12484
rect 19992 12540 20056 12544
rect 19992 12484 19996 12540
rect 19996 12484 20052 12540
rect 20052 12484 20056 12540
rect 19992 12480 20056 12484
rect 20072 12540 20136 12544
rect 20072 12484 20076 12540
rect 20076 12484 20132 12540
rect 20132 12484 20136 12540
rect 20072 12480 20136 12484
rect 20152 12540 20216 12544
rect 20152 12484 20156 12540
rect 20156 12484 20212 12540
rect 20212 12484 20216 12540
rect 20152 12480 20216 12484
rect 20232 12540 20296 12544
rect 20232 12484 20236 12540
rect 20236 12484 20292 12540
rect 20292 12484 20296 12540
rect 20232 12480 20296 12484
rect 2652 11996 2716 12000
rect 2652 11940 2656 11996
rect 2656 11940 2712 11996
rect 2712 11940 2716 11996
rect 2652 11936 2716 11940
rect 2732 11996 2796 12000
rect 2732 11940 2736 11996
rect 2736 11940 2792 11996
rect 2792 11940 2796 11996
rect 2732 11936 2796 11940
rect 2812 11996 2876 12000
rect 2812 11940 2816 11996
rect 2816 11940 2872 11996
rect 2872 11940 2876 11996
rect 2812 11936 2876 11940
rect 2892 11996 2956 12000
rect 2892 11940 2896 11996
rect 2896 11940 2952 11996
rect 2952 11940 2956 11996
rect 2892 11936 2956 11940
rect 2972 11996 3036 12000
rect 2972 11940 2976 11996
rect 2976 11940 3032 11996
rect 3032 11940 3036 11996
rect 2972 11936 3036 11940
rect 8652 11996 8716 12000
rect 8652 11940 8656 11996
rect 8656 11940 8712 11996
rect 8712 11940 8716 11996
rect 8652 11936 8716 11940
rect 8732 11996 8796 12000
rect 8732 11940 8736 11996
rect 8736 11940 8792 11996
rect 8792 11940 8796 11996
rect 8732 11936 8796 11940
rect 8812 11996 8876 12000
rect 8812 11940 8816 11996
rect 8816 11940 8872 11996
rect 8872 11940 8876 11996
rect 8812 11936 8876 11940
rect 8892 11996 8956 12000
rect 8892 11940 8896 11996
rect 8896 11940 8952 11996
rect 8952 11940 8956 11996
rect 8892 11936 8956 11940
rect 8972 11996 9036 12000
rect 8972 11940 8976 11996
rect 8976 11940 9032 11996
rect 9032 11940 9036 11996
rect 8972 11936 9036 11940
rect 14652 11996 14716 12000
rect 14652 11940 14656 11996
rect 14656 11940 14712 11996
rect 14712 11940 14716 11996
rect 14652 11936 14716 11940
rect 14732 11996 14796 12000
rect 14732 11940 14736 11996
rect 14736 11940 14792 11996
rect 14792 11940 14796 11996
rect 14732 11936 14796 11940
rect 14812 11996 14876 12000
rect 14812 11940 14816 11996
rect 14816 11940 14872 11996
rect 14872 11940 14876 11996
rect 14812 11936 14876 11940
rect 14892 11996 14956 12000
rect 14892 11940 14896 11996
rect 14896 11940 14952 11996
rect 14952 11940 14956 11996
rect 14892 11936 14956 11940
rect 14972 11996 15036 12000
rect 14972 11940 14976 11996
rect 14976 11940 15032 11996
rect 15032 11940 15036 11996
rect 14972 11936 15036 11940
rect 20652 11996 20716 12000
rect 20652 11940 20656 11996
rect 20656 11940 20712 11996
rect 20712 11940 20716 11996
rect 20652 11936 20716 11940
rect 20732 11996 20796 12000
rect 20732 11940 20736 11996
rect 20736 11940 20792 11996
rect 20792 11940 20796 11996
rect 20732 11936 20796 11940
rect 20812 11996 20876 12000
rect 20812 11940 20816 11996
rect 20816 11940 20872 11996
rect 20872 11940 20876 11996
rect 20812 11936 20876 11940
rect 20892 11996 20956 12000
rect 20892 11940 20896 11996
rect 20896 11940 20952 11996
rect 20952 11940 20956 11996
rect 20892 11936 20956 11940
rect 20972 11996 21036 12000
rect 20972 11940 20976 11996
rect 20976 11940 21032 11996
rect 21032 11940 21036 11996
rect 20972 11936 21036 11940
rect 1912 11452 1976 11456
rect 1912 11396 1916 11452
rect 1916 11396 1972 11452
rect 1972 11396 1976 11452
rect 1912 11392 1976 11396
rect 1992 11452 2056 11456
rect 1992 11396 1996 11452
rect 1996 11396 2052 11452
rect 2052 11396 2056 11452
rect 1992 11392 2056 11396
rect 2072 11452 2136 11456
rect 2072 11396 2076 11452
rect 2076 11396 2132 11452
rect 2132 11396 2136 11452
rect 2072 11392 2136 11396
rect 2152 11452 2216 11456
rect 2152 11396 2156 11452
rect 2156 11396 2212 11452
rect 2212 11396 2216 11452
rect 2152 11392 2216 11396
rect 2232 11452 2296 11456
rect 2232 11396 2236 11452
rect 2236 11396 2292 11452
rect 2292 11396 2296 11452
rect 2232 11392 2296 11396
rect 7912 11452 7976 11456
rect 7912 11396 7916 11452
rect 7916 11396 7972 11452
rect 7972 11396 7976 11452
rect 7912 11392 7976 11396
rect 7992 11452 8056 11456
rect 7992 11396 7996 11452
rect 7996 11396 8052 11452
rect 8052 11396 8056 11452
rect 7992 11392 8056 11396
rect 8072 11452 8136 11456
rect 8072 11396 8076 11452
rect 8076 11396 8132 11452
rect 8132 11396 8136 11452
rect 8072 11392 8136 11396
rect 8152 11452 8216 11456
rect 8152 11396 8156 11452
rect 8156 11396 8212 11452
rect 8212 11396 8216 11452
rect 8152 11392 8216 11396
rect 8232 11452 8296 11456
rect 8232 11396 8236 11452
rect 8236 11396 8292 11452
rect 8292 11396 8296 11452
rect 8232 11392 8296 11396
rect 13912 11452 13976 11456
rect 13912 11396 13916 11452
rect 13916 11396 13972 11452
rect 13972 11396 13976 11452
rect 13912 11392 13976 11396
rect 13992 11452 14056 11456
rect 13992 11396 13996 11452
rect 13996 11396 14052 11452
rect 14052 11396 14056 11452
rect 13992 11392 14056 11396
rect 14072 11452 14136 11456
rect 14072 11396 14076 11452
rect 14076 11396 14132 11452
rect 14132 11396 14136 11452
rect 14072 11392 14136 11396
rect 14152 11452 14216 11456
rect 14152 11396 14156 11452
rect 14156 11396 14212 11452
rect 14212 11396 14216 11452
rect 14152 11392 14216 11396
rect 14232 11452 14296 11456
rect 14232 11396 14236 11452
rect 14236 11396 14292 11452
rect 14292 11396 14296 11452
rect 14232 11392 14296 11396
rect 19912 11452 19976 11456
rect 19912 11396 19916 11452
rect 19916 11396 19972 11452
rect 19972 11396 19976 11452
rect 19912 11392 19976 11396
rect 19992 11452 20056 11456
rect 19992 11396 19996 11452
rect 19996 11396 20052 11452
rect 20052 11396 20056 11452
rect 19992 11392 20056 11396
rect 20072 11452 20136 11456
rect 20072 11396 20076 11452
rect 20076 11396 20132 11452
rect 20132 11396 20136 11452
rect 20072 11392 20136 11396
rect 20152 11452 20216 11456
rect 20152 11396 20156 11452
rect 20156 11396 20212 11452
rect 20212 11396 20216 11452
rect 20152 11392 20216 11396
rect 20232 11452 20296 11456
rect 20232 11396 20236 11452
rect 20236 11396 20292 11452
rect 20292 11396 20296 11452
rect 20232 11392 20296 11396
rect 2652 10908 2716 10912
rect 2652 10852 2656 10908
rect 2656 10852 2712 10908
rect 2712 10852 2716 10908
rect 2652 10848 2716 10852
rect 2732 10908 2796 10912
rect 2732 10852 2736 10908
rect 2736 10852 2792 10908
rect 2792 10852 2796 10908
rect 2732 10848 2796 10852
rect 2812 10908 2876 10912
rect 2812 10852 2816 10908
rect 2816 10852 2872 10908
rect 2872 10852 2876 10908
rect 2812 10848 2876 10852
rect 2892 10908 2956 10912
rect 2892 10852 2896 10908
rect 2896 10852 2952 10908
rect 2952 10852 2956 10908
rect 2892 10848 2956 10852
rect 2972 10908 3036 10912
rect 2972 10852 2976 10908
rect 2976 10852 3032 10908
rect 3032 10852 3036 10908
rect 2972 10848 3036 10852
rect 8652 10908 8716 10912
rect 8652 10852 8656 10908
rect 8656 10852 8712 10908
rect 8712 10852 8716 10908
rect 8652 10848 8716 10852
rect 8732 10908 8796 10912
rect 8732 10852 8736 10908
rect 8736 10852 8792 10908
rect 8792 10852 8796 10908
rect 8732 10848 8796 10852
rect 8812 10908 8876 10912
rect 8812 10852 8816 10908
rect 8816 10852 8872 10908
rect 8872 10852 8876 10908
rect 8812 10848 8876 10852
rect 8892 10908 8956 10912
rect 8892 10852 8896 10908
rect 8896 10852 8952 10908
rect 8952 10852 8956 10908
rect 8892 10848 8956 10852
rect 8972 10908 9036 10912
rect 8972 10852 8976 10908
rect 8976 10852 9032 10908
rect 9032 10852 9036 10908
rect 8972 10848 9036 10852
rect 14652 10908 14716 10912
rect 14652 10852 14656 10908
rect 14656 10852 14712 10908
rect 14712 10852 14716 10908
rect 14652 10848 14716 10852
rect 14732 10908 14796 10912
rect 14732 10852 14736 10908
rect 14736 10852 14792 10908
rect 14792 10852 14796 10908
rect 14732 10848 14796 10852
rect 14812 10908 14876 10912
rect 14812 10852 14816 10908
rect 14816 10852 14872 10908
rect 14872 10852 14876 10908
rect 14812 10848 14876 10852
rect 14892 10908 14956 10912
rect 14892 10852 14896 10908
rect 14896 10852 14952 10908
rect 14952 10852 14956 10908
rect 14892 10848 14956 10852
rect 14972 10908 15036 10912
rect 14972 10852 14976 10908
rect 14976 10852 15032 10908
rect 15032 10852 15036 10908
rect 14972 10848 15036 10852
rect 20652 10908 20716 10912
rect 20652 10852 20656 10908
rect 20656 10852 20712 10908
rect 20712 10852 20716 10908
rect 20652 10848 20716 10852
rect 20732 10908 20796 10912
rect 20732 10852 20736 10908
rect 20736 10852 20792 10908
rect 20792 10852 20796 10908
rect 20732 10848 20796 10852
rect 20812 10908 20876 10912
rect 20812 10852 20816 10908
rect 20816 10852 20872 10908
rect 20872 10852 20876 10908
rect 20812 10848 20876 10852
rect 20892 10908 20956 10912
rect 20892 10852 20896 10908
rect 20896 10852 20952 10908
rect 20952 10852 20956 10908
rect 20892 10848 20956 10852
rect 20972 10908 21036 10912
rect 20972 10852 20976 10908
rect 20976 10852 21032 10908
rect 21032 10852 21036 10908
rect 20972 10848 21036 10852
rect 9444 10644 9508 10708
rect 1912 10364 1976 10368
rect 1912 10308 1916 10364
rect 1916 10308 1972 10364
rect 1972 10308 1976 10364
rect 1912 10304 1976 10308
rect 1992 10364 2056 10368
rect 1992 10308 1996 10364
rect 1996 10308 2052 10364
rect 2052 10308 2056 10364
rect 1992 10304 2056 10308
rect 2072 10364 2136 10368
rect 2072 10308 2076 10364
rect 2076 10308 2132 10364
rect 2132 10308 2136 10364
rect 2072 10304 2136 10308
rect 2152 10364 2216 10368
rect 2152 10308 2156 10364
rect 2156 10308 2212 10364
rect 2212 10308 2216 10364
rect 2152 10304 2216 10308
rect 2232 10364 2296 10368
rect 2232 10308 2236 10364
rect 2236 10308 2292 10364
rect 2292 10308 2296 10364
rect 2232 10304 2296 10308
rect 7912 10364 7976 10368
rect 7912 10308 7916 10364
rect 7916 10308 7972 10364
rect 7972 10308 7976 10364
rect 7912 10304 7976 10308
rect 7992 10364 8056 10368
rect 7992 10308 7996 10364
rect 7996 10308 8052 10364
rect 8052 10308 8056 10364
rect 7992 10304 8056 10308
rect 8072 10364 8136 10368
rect 8072 10308 8076 10364
rect 8076 10308 8132 10364
rect 8132 10308 8136 10364
rect 8072 10304 8136 10308
rect 8152 10364 8216 10368
rect 8152 10308 8156 10364
rect 8156 10308 8212 10364
rect 8212 10308 8216 10364
rect 8152 10304 8216 10308
rect 8232 10364 8296 10368
rect 8232 10308 8236 10364
rect 8236 10308 8292 10364
rect 8292 10308 8296 10364
rect 8232 10304 8296 10308
rect 13912 10364 13976 10368
rect 13912 10308 13916 10364
rect 13916 10308 13972 10364
rect 13972 10308 13976 10364
rect 13912 10304 13976 10308
rect 13992 10364 14056 10368
rect 13992 10308 13996 10364
rect 13996 10308 14052 10364
rect 14052 10308 14056 10364
rect 13992 10304 14056 10308
rect 14072 10364 14136 10368
rect 14072 10308 14076 10364
rect 14076 10308 14132 10364
rect 14132 10308 14136 10364
rect 14072 10304 14136 10308
rect 14152 10364 14216 10368
rect 14152 10308 14156 10364
rect 14156 10308 14212 10364
rect 14212 10308 14216 10364
rect 14152 10304 14216 10308
rect 14232 10364 14296 10368
rect 14232 10308 14236 10364
rect 14236 10308 14292 10364
rect 14292 10308 14296 10364
rect 14232 10304 14296 10308
rect 19912 10364 19976 10368
rect 19912 10308 19916 10364
rect 19916 10308 19972 10364
rect 19972 10308 19976 10364
rect 19912 10304 19976 10308
rect 19992 10364 20056 10368
rect 19992 10308 19996 10364
rect 19996 10308 20052 10364
rect 20052 10308 20056 10364
rect 19992 10304 20056 10308
rect 20072 10364 20136 10368
rect 20072 10308 20076 10364
rect 20076 10308 20132 10364
rect 20132 10308 20136 10364
rect 20072 10304 20136 10308
rect 20152 10364 20216 10368
rect 20152 10308 20156 10364
rect 20156 10308 20212 10364
rect 20212 10308 20216 10364
rect 20152 10304 20216 10308
rect 20232 10364 20296 10368
rect 20232 10308 20236 10364
rect 20236 10308 20292 10364
rect 20292 10308 20296 10364
rect 20232 10304 20296 10308
rect 2652 9820 2716 9824
rect 2652 9764 2656 9820
rect 2656 9764 2712 9820
rect 2712 9764 2716 9820
rect 2652 9760 2716 9764
rect 2732 9820 2796 9824
rect 2732 9764 2736 9820
rect 2736 9764 2792 9820
rect 2792 9764 2796 9820
rect 2732 9760 2796 9764
rect 2812 9820 2876 9824
rect 2812 9764 2816 9820
rect 2816 9764 2872 9820
rect 2872 9764 2876 9820
rect 2812 9760 2876 9764
rect 2892 9820 2956 9824
rect 2892 9764 2896 9820
rect 2896 9764 2952 9820
rect 2952 9764 2956 9820
rect 2892 9760 2956 9764
rect 2972 9820 3036 9824
rect 2972 9764 2976 9820
rect 2976 9764 3032 9820
rect 3032 9764 3036 9820
rect 2972 9760 3036 9764
rect 8652 9820 8716 9824
rect 8652 9764 8656 9820
rect 8656 9764 8712 9820
rect 8712 9764 8716 9820
rect 8652 9760 8716 9764
rect 8732 9820 8796 9824
rect 8732 9764 8736 9820
rect 8736 9764 8792 9820
rect 8792 9764 8796 9820
rect 8732 9760 8796 9764
rect 8812 9820 8876 9824
rect 8812 9764 8816 9820
rect 8816 9764 8872 9820
rect 8872 9764 8876 9820
rect 8812 9760 8876 9764
rect 8892 9820 8956 9824
rect 8892 9764 8896 9820
rect 8896 9764 8952 9820
rect 8952 9764 8956 9820
rect 8892 9760 8956 9764
rect 8972 9820 9036 9824
rect 8972 9764 8976 9820
rect 8976 9764 9032 9820
rect 9032 9764 9036 9820
rect 8972 9760 9036 9764
rect 14652 9820 14716 9824
rect 14652 9764 14656 9820
rect 14656 9764 14712 9820
rect 14712 9764 14716 9820
rect 14652 9760 14716 9764
rect 14732 9820 14796 9824
rect 14732 9764 14736 9820
rect 14736 9764 14792 9820
rect 14792 9764 14796 9820
rect 14732 9760 14796 9764
rect 14812 9820 14876 9824
rect 14812 9764 14816 9820
rect 14816 9764 14872 9820
rect 14872 9764 14876 9820
rect 14812 9760 14876 9764
rect 14892 9820 14956 9824
rect 14892 9764 14896 9820
rect 14896 9764 14952 9820
rect 14952 9764 14956 9820
rect 14892 9760 14956 9764
rect 14972 9820 15036 9824
rect 14972 9764 14976 9820
rect 14976 9764 15032 9820
rect 15032 9764 15036 9820
rect 14972 9760 15036 9764
rect 20652 9820 20716 9824
rect 20652 9764 20656 9820
rect 20656 9764 20712 9820
rect 20712 9764 20716 9820
rect 20652 9760 20716 9764
rect 20732 9820 20796 9824
rect 20732 9764 20736 9820
rect 20736 9764 20792 9820
rect 20792 9764 20796 9820
rect 20732 9760 20796 9764
rect 20812 9820 20876 9824
rect 20812 9764 20816 9820
rect 20816 9764 20872 9820
rect 20872 9764 20876 9820
rect 20812 9760 20876 9764
rect 20892 9820 20956 9824
rect 20892 9764 20896 9820
rect 20896 9764 20952 9820
rect 20952 9764 20956 9820
rect 20892 9760 20956 9764
rect 20972 9820 21036 9824
rect 20972 9764 20976 9820
rect 20976 9764 21032 9820
rect 21032 9764 21036 9820
rect 20972 9760 21036 9764
rect 1912 9276 1976 9280
rect 1912 9220 1916 9276
rect 1916 9220 1972 9276
rect 1972 9220 1976 9276
rect 1912 9216 1976 9220
rect 1992 9276 2056 9280
rect 1992 9220 1996 9276
rect 1996 9220 2052 9276
rect 2052 9220 2056 9276
rect 1992 9216 2056 9220
rect 2072 9276 2136 9280
rect 2072 9220 2076 9276
rect 2076 9220 2132 9276
rect 2132 9220 2136 9276
rect 2072 9216 2136 9220
rect 2152 9276 2216 9280
rect 2152 9220 2156 9276
rect 2156 9220 2212 9276
rect 2212 9220 2216 9276
rect 2152 9216 2216 9220
rect 2232 9276 2296 9280
rect 2232 9220 2236 9276
rect 2236 9220 2292 9276
rect 2292 9220 2296 9276
rect 2232 9216 2296 9220
rect 7912 9276 7976 9280
rect 7912 9220 7916 9276
rect 7916 9220 7972 9276
rect 7972 9220 7976 9276
rect 7912 9216 7976 9220
rect 7992 9276 8056 9280
rect 7992 9220 7996 9276
rect 7996 9220 8052 9276
rect 8052 9220 8056 9276
rect 7992 9216 8056 9220
rect 8072 9276 8136 9280
rect 8072 9220 8076 9276
rect 8076 9220 8132 9276
rect 8132 9220 8136 9276
rect 8072 9216 8136 9220
rect 8152 9276 8216 9280
rect 8152 9220 8156 9276
rect 8156 9220 8212 9276
rect 8212 9220 8216 9276
rect 8152 9216 8216 9220
rect 8232 9276 8296 9280
rect 8232 9220 8236 9276
rect 8236 9220 8292 9276
rect 8292 9220 8296 9276
rect 8232 9216 8296 9220
rect 13912 9276 13976 9280
rect 13912 9220 13916 9276
rect 13916 9220 13972 9276
rect 13972 9220 13976 9276
rect 13912 9216 13976 9220
rect 13992 9276 14056 9280
rect 13992 9220 13996 9276
rect 13996 9220 14052 9276
rect 14052 9220 14056 9276
rect 13992 9216 14056 9220
rect 14072 9276 14136 9280
rect 14072 9220 14076 9276
rect 14076 9220 14132 9276
rect 14132 9220 14136 9276
rect 14072 9216 14136 9220
rect 14152 9276 14216 9280
rect 14152 9220 14156 9276
rect 14156 9220 14212 9276
rect 14212 9220 14216 9276
rect 14152 9216 14216 9220
rect 14232 9276 14296 9280
rect 14232 9220 14236 9276
rect 14236 9220 14292 9276
rect 14292 9220 14296 9276
rect 14232 9216 14296 9220
rect 19912 9276 19976 9280
rect 19912 9220 19916 9276
rect 19916 9220 19972 9276
rect 19972 9220 19976 9276
rect 19912 9216 19976 9220
rect 19992 9276 20056 9280
rect 19992 9220 19996 9276
rect 19996 9220 20052 9276
rect 20052 9220 20056 9276
rect 19992 9216 20056 9220
rect 20072 9276 20136 9280
rect 20072 9220 20076 9276
rect 20076 9220 20132 9276
rect 20132 9220 20136 9276
rect 20072 9216 20136 9220
rect 20152 9276 20216 9280
rect 20152 9220 20156 9276
rect 20156 9220 20212 9276
rect 20212 9220 20216 9276
rect 20152 9216 20216 9220
rect 20232 9276 20296 9280
rect 20232 9220 20236 9276
rect 20236 9220 20292 9276
rect 20292 9220 20296 9276
rect 20232 9216 20296 9220
rect 2652 8732 2716 8736
rect 2652 8676 2656 8732
rect 2656 8676 2712 8732
rect 2712 8676 2716 8732
rect 2652 8672 2716 8676
rect 2732 8732 2796 8736
rect 2732 8676 2736 8732
rect 2736 8676 2792 8732
rect 2792 8676 2796 8732
rect 2732 8672 2796 8676
rect 2812 8732 2876 8736
rect 2812 8676 2816 8732
rect 2816 8676 2872 8732
rect 2872 8676 2876 8732
rect 2812 8672 2876 8676
rect 2892 8732 2956 8736
rect 2892 8676 2896 8732
rect 2896 8676 2952 8732
rect 2952 8676 2956 8732
rect 2892 8672 2956 8676
rect 2972 8732 3036 8736
rect 2972 8676 2976 8732
rect 2976 8676 3032 8732
rect 3032 8676 3036 8732
rect 2972 8672 3036 8676
rect 8652 8732 8716 8736
rect 8652 8676 8656 8732
rect 8656 8676 8712 8732
rect 8712 8676 8716 8732
rect 8652 8672 8716 8676
rect 8732 8732 8796 8736
rect 8732 8676 8736 8732
rect 8736 8676 8792 8732
rect 8792 8676 8796 8732
rect 8732 8672 8796 8676
rect 8812 8732 8876 8736
rect 8812 8676 8816 8732
rect 8816 8676 8872 8732
rect 8872 8676 8876 8732
rect 8812 8672 8876 8676
rect 8892 8732 8956 8736
rect 8892 8676 8896 8732
rect 8896 8676 8952 8732
rect 8952 8676 8956 8732
rect 8892 8672 8956 8676
rect 8972 8732 9036 8736
rect 8972 8676 8976 8732
rect 8976 8676 9032 8732
rect 9032 8676 9036 8732
rect 8972 8672 9036 8676
rect 14652 8732 14716 8736
rect 14652 8676 14656 8732
rect 14656 8676 14712 8732
rect 14712 8676 14716 8732
rect 14652 8672 14716 8676
rect 14732 8732 14796 8736
rect 14732 8676 14736 8732
rect 14736 8676 14792 8732
rect 14792 8676 14796 8732
rect 14732 8672 14796 8676
rect 14812 8732 14876 8736
rect 14812 8676 14816 8732
rect 14816 8676 14872 8732
rect 14872 8676 14876 8732
rect 14812 8672 14876 8676
rect 14892 8732 14956 8736
rect 14892 8676 14896 8732
rect 14896 8676 14952 8732
rect 14952 8676 14956 8732
rect 14892 8672 14956 8676
rect 14972 8732 15036 8736
rect 14972 8676 14976 8732
rect 14976 8676 15032 8732
rect 15032 8676 15036 8732
rect 14972 8672 15036 8676
rect 20652 8732 20716 8736
rect 20652 8676 20656 8732
rect 20656 8676 20712 8732
rect 20712 8676 20716 8732
rect 20652 8672 20716 8676
rect 20732 8732 20796 8736
rect 20732 8676 20736 8732
rect 20736 8676 20792 8732
rect 20792 8676 20796 8732
rect 20732 8672 20796 8676
rect 20812 8732 20876 8736
rect 20812 8676 20816 8732
rect 20816 8676 20872 8732
rect 20872 8676 20876 8732
rect 20812 8672 20876 8676
rect 20892 8732 20956 8736
rect 20892 8676 20896 8732
rect 20896 8676 20952 8732
rect 20952 8676 20956 8732
rect 20892 8672 20956 8676
rect 20972 8732 21036 8736
rect 20972 8676 20976 8732
rect 20976 8676 21032 8732
rect 21032 8676 21036 8732
rect 20972 8672 21036 8676
rect 1912 8188 1976 8192
rect 1912 8132 1916 8188
rect 1916 8132 1972 8188
rect 1972 8132 1976 8188
rect 1912 8128 1976 8132
rect 1992 8188 2056 8192
rect 1992 8132 1996 8188
rect 1996 8132 2052 8188
rect 2052 8132 2056 8188
rect 1992 8128 2056 8132
rect 2072 8188 2136 8192
rect 2072 8132 2076 8188
rect 2076 8132 2132 8188
rect 2132 8132 2136 8188
rect 2072 8128 2136 8132
rect 2152 8188 2216 8192
rect 2152 8132 2156 8188
rect 2156 8132 2212 8188
rect 2212 8132 2216 8188
rect 2152 8128 2216 8132
rect 2232 8188 2296 8192
rect 2232 8132 2236 8188
rect 2236 8132 2292 8188
rect 2292 8132 2296 8188
rect 2232 8128 2296 8132
rect 7912 8188 7976 8192
rect 7912 8132 7916 8188
rect 7916 8132 7972 8188
rect 7972 8132 7976 8188
rect 7912 8128 7976 8132
rect 7992 8188 8056 8192
rect 7992 8132 7996 8188
rect 7996 8132 8052 8188
rect 8052 8132 8056 8188
rect 7992 8128 8056 8132
rect 8072 8188 8136 8192
rect 8072 8132 8076 8188
rect 8076 8132 8132 8188
rect 8132 8132 8136 8188
rect 8072 8128 8136 8132
rect 8152 8188 8216 8192
rect 8152 8132 8156 8188
rect 8156 8132 8212 8188
rect 8212 8132 8216 8188
rect 8152 8128 8216 8132
rect 8232 8188 8296 8192
rect 8232 8132 8236 8188
rect 8236 8132 8292 8188
rect 8292 8132 8296 8188
rect 8232 8128 8296 8132
rect 13912 8188 13976 8192
rect 13912 8132 13916 8188
rect 13916 8132 13972 8188
rect 13972 8132 13976 8188
rect 13912 8128 13976 8132
rect 13992 8188 14056 8192
rect 13992 8132 13996 8188
rect 13996 8132 14052 8188
rect 14052 8132 14056 8188
rect 13992 8128 14056 8132
rect 14072 8188 14136 8192
rect 14072 8132 14076 8188
rect 14076 8132 14132 8188
rect 14132 8132 14136 8188
rect 14072 8128 14136 8132
rect 14152 8188 14216 8192
rect 14152 8132 14156 8188
rect 14156 8132 14212 8188
rect 14212 8132 14216 8188
rect 14152 8128 14216 8132
rect 14232 8188 14296 8192
rect 14232 8132 14236 8188
rect 14236 8132 14292 8188
rect 14292 8132 14296 8188
rect 14232 8128 14296 8132
rect 19912 8188 19976 8192
rect 19912 8132 19916 8188
rect 19916 8132 19972 8188
rect 19972 8132 19976 8188
rect 19912 8128 19976 8132
rect 19992 8188 20056 8192
rect 19992 8132 19996 8188
rect 19996 8132 20052 8188
rect 20052 8132 20056 8188
rect 19992 8128 20056 8132
rect 20072 8188 20136 8192
rect 20072 8132 20076 8188
rect 20076 8132 20132 8188
rect 20132 8132 20136 8188
rect 20072 8128 20136 8132
rect 20152 8188 20216 8192
rect 20152 8132 20156 8188
rect 20156 8132 20212 8188
rect 20212 8132 20216 8188
rect 20152 8128 20216 8132
rect 20232 8188 20296 8192
rect 20232 8132 20236 8188
rect 20236 8132 20292 8188
rect 20292 8132 20296 8188
rect 20232 8128 20296 8132
rect 2652 7644 2716 7648
rect 2652 7588 2656 7644
rect 2656 7588 2712 7644
rect 2712 7588 2716 7644
rect 2652 7584 2716 7588
rect 2732 7644 2796 7648
rect 2732 7588 2736 7644
rect 2736 7588 2792 7644
rect 2792 7588 2796 7644
rect 2732 7584 2796 7588
rect 2812 7644 2876 7648
rect 2812 7588 2816 7644
rect 2816 7588 2872 7644
rect 2872 7588 2876 7644
rect 2812 7584 2876 7588
rect 2892 7644 2956 7648
rect 2892 7588 2896 7644
rect 2896 7588 2952 7644
rect 2952 7588 2956 7644
rect 2892 7584 2956 7588
rect 2972 7644 3036 7648
rect 2972 7588 2976 7644
rect 2976 7588 3032 7644
rect 3032 7588 3036 7644
rect 2972 7584 3036 7588
rect 8652 7644 8716 7648
rect 8652 7588 8656 7644
rect 8656 7588 8712 7644
rect 8712 7588 8716 7644
rect 8652 7584 8716 7588
rect 8732 7644 8796 7648
rect 8732 7588 8736 7644
rect 8736 7588 8792 7644
rect 8792 7588 8796 7644
rect 8732 7584 8796 7588
rect 8812 7644 8876 7648
rect 8812 7588 8816 7644
rect 8816 7588 8872 7644
rect 8872 7588 8876 7644
rect 8812 7584 8876 7588
rect 8892 7644 8956 7648
rect 8892 7588 8896 7644
rect 8896 7588 8952 7644
rect 8952 7588 8956 7644
rect 8892 7584 8956 7588
rect 8972 7644 9036 7648
rect 8972 7588 8976 7644
rect 8976 7588 9032 7644
rect 9032 7588 9036 7644
rect 8972 7584 9036 7588
rect 14652 7644 14716 7648
rect 14652 7588 14656 7644
rect 14656 7588 14712 7644
rect 14712 7588 14716 7644
rect 14652 7584 14716 7588
rect 14732 7644 14796 7648
rect 14732 7588 14736 7644
rect 14736 7588 14792 7644
rect 14792 7588 14796 7644
rect 14732 7584 14796 7588
rect 14812 7644 14876 7648
rect 14812 7588 14816 7644
rect 14816 7588 14872 7644
rect 14872 7588 14876 7644
rect 14812 7584 14876 7588
rect 14892 7644 14956 7648
rect 14892 7588 14896 7644
rect 14896 7588 14952 7644
rect 14952 7588 14956 7644
rect 14892 7584 14956 7588
rect 14972 7644 15036 7648
rect 14972 7588 14976 7644
rect 14976 7588 15032 7644
rect 15032 7588 15036 7644
rect 14972 7584 15036 7588
rect 20652 7644 20716 7648
rect 20652 7588 20656 7644
rect 20656 7588 20712 7644
rect 20712 7588 20716 7644
rect 20652 7584 20716 7588
rect 20732 7644 20796 7648
rect 20732 7588 20736 7644
rect 20736 7588 20792 7644
rect 20792 7588 20796 7644
rect 20732 7584 20796 7588
rect 20812 7644 20876 7648
rect 20812 7588 20816 7644
rect 20816 7588 20872 7644
rect 20872 7588 20876 7644
rect 20812 7584 20876 7588
rect 20892 7644 20956 7648
rect 20892 7588 20896 7644
rect 20896 7588 20952 7644
rect 20952 7588 20956 7644
rect 20892 7584 20956 7588
rect 20972 7644 21036 7648
rect 20972 7588 20976 7644
rect 20976 7588 21032 7644
rect 21032 7588 21036 7644
rect 20972 7584 21036 7588
rect 1912 7100 1976 7104
rect 1912 7044 1916 7100
rect 1916 7044 1972 7100
rect 1972 7044 1976 7100
rect 1912 7040 1976 7044
rect 1992 7100 2056 7104
rect 1992 7044 1996 7100
rect 1996 7044 2052 7100
rect 2052 7044 2056 7100
rect 1992 7040 2056 7044
rect 2072 7100 2136 7104
rect 2072 7044 2076 7100
rect 2076 7044 2132 7100
rect 2132 7044 2136 7100
rect 2072 7040 2136 7044
rect 2152 7100 2216 7104
rect 2152 7044 2156 7100
rect 2156 7044 2212 7100
rect 2212 7044 2216 7100
rect 2152 7040 2216 7044
rect 2232 7100 2296 7104
rect 2232 7044 2236 7100
rect 2236 7044 2292 7100
rect 2292 7044 2296 7100
rect 2232 7040 2296 7044
rect 7912 7100 7976 7104
rect 7912 7044 7916 7100
rect 7916 7044 7972 7100
rect 7972 7044 7976 7100
rect 7912 7040 7976 7044
rect 7992 7100 8056 7104
rect 7992 7044 7996 7100
rect 7996 7044 8052 7100
rect 8052 7044 8056 7100
rect 7992 7040 8056 7044
rect 8072 7100 8136 7104
rect 8072 7044 8076 7100
rect 8076 7044 8132 7100
rect 8132 7044 8136 7100
rect 8072 7040 8136 7044
rect 8152 7100 8216 7104
rect 8152 7044 8156 7100
rect 8156 7044 8212 7100
rect 8212 7044 8216 7100
rect 8152 7040 8216 7044
rect 8232 7100 8296 7104
rect 8232 7044 8236 7100
rect 8236 7044 8292 7100
rect 8292 7044 8296 7100
rect 8232 7040 8296 7044
rect 13912 7100 13976 7104
rect 13912 7044 13916 7100
rect 13916 7044 13972 7100
rect 13972 7044 13976 7100
rect 13912 7040 13976 7044
rect 13992 7100 14056 7104
rect 13992 7044 13996 7100
rect 13996 7044 14052 7100
rect 14052 7044 14056 7100
rect 13992 7040 14056 7044
rect 14072 7100 14136 7104
rect 14072 7044 14076 7100
rect 14076 7044 14132 7100
rect 14132 7044 14136 7100
rect 14072 7040 14136 7044
rect 14152 7100 14216 7104
rect 14152 7044 14156 7100
rect 14156 7044 14212 7100
rect 14212 7044 14216 7100
rect 14152 7040 14216 7044
rect 14232 7100 14296 7104
rect 14232 7044 14236 7100
rect 14236 7044 14292 7100
rect 14292 7044 14296 7100
rect 14232 7040 14296 7044
rect 19912 7100 19976 7104
rect 19912 7044 19916 7100
rect 19916 7044 19972 7100
rect 19972 7044 19976 7100
rect 19912 7040 19976 7044
rect 19992 7100 20056 7104
rect 19992 7044 19996 7100
rect 19996 7044 20052 7100
rect 20052 7044 20056 7100
rect 19992 7040 20056 7044
rect 20072 7100 20136 7104
rect 20072 7044 20076 7100
rect 20076 7044 20132 7100
rect 20132 7044 20136 7100
rect 20072 7040 20136 7044
rect 20152 7100 20216 7104
rect 20152 7044 20156 7100
rect 20156 7044 20212 7100
rect 20212 7044 20216 7100
rect 20152 7040 20216 7044
rect 20232 7100 20296 7104
rect 20232 7044 20236 7100
rect 20236 7044 20292 7100
rect 20292 7044 20296 7100
rect 20232 7040 20296 7044
rect 2652 6556 2716 6560
rect 2652 6500 2656 6556
rect 2656 6500 2712 6556
rect 2712 6500 2716 6556
rect 2652 6496 2716 6500
rect 2732 6556 2796 6560
rect 2732 6500 2736 6556
rect 2736 6500 2792 6556
rect 2792 6500 2796 6556
rect 2732 6496 2796 6500
rect 2812 6556 2876 6560
rect 2812 6500 2816 6556
rect 2816 6500 2872 6556
rect 2872 6500 2876 6556
rect 2812 6496 2876 6500
rect 2892 6556 2956 6560
rect 2892 6500 2896 6556
rect 2896 6500 2952 6556
rect 2952 6500 2956 6556
rect 2892 6496 2956 6500
rect 2972 6556 3036 6560
rect 2972 6500 2976 6556
rect 2976 6500 3032 6556
rect 3032 6500 3036 6556
rect 2972 6496 3036 6500
rect 8652 6556 8716 6560
rect 8652 6500 8656 6556
rect 8656 6500 8712 6556
rect 8712 6500 8716 6556
rect 8652 6496 8716 6500
rect 8732 6556 8796 6560
rect 8732 6500 8736 6556
rect 8736 6500 8792 6556
rect 8792 6500 8796 6556
rect 8732 6496 8796 6500
rect 8812 6556 8876 6560
rect 8812 6500 8816 6556
rect 8816 6500 8872 6556
rect 8872 6500 8876 6556
rect 8812 6496 8876 6500
rect 8892 6556 8956 6560
rect 8892 6500 8896 6556
rect 8896 6500 8952 6556
rect 8952 6500 8956 6556
rect 8892 6496 8956 6500
rect 8972 6556 9036 6560
rect 8972 6500 8976 6556
rect 8976 6500 9032 6556
rect 9032 6500 9036 6556
rect 8972 6496 9036 6500
rect 14652 6556 14716 6560
rect 14652 6500 14656 6556
rect 14656 6500 14712 6556
rect 14712 6500 14716 6556
rect 14652 6496 14716 6500
rect 14732 6556 14796 6560
rect 14732 6500 14736 6556
rect 14736 6500 14792 6556
rect 14792 6500 14796 6556
rect 14732 6496 14796 6500
rect 14812 6556 14876 6560
rect 14812 6500 14816 6556
rect 14816 6500 14872 6556
rect 14872 6500 14876 6556
rect 14812 6496 14876 6500
rect 14892 6556 14956 6560
rect 14892 6500 14896 6556
rect 14896 6500 14952 6556
rect 14952 6500 14956 6556
rect 14892 6496 14956 6500
rect 14972 6556 15036 6560
rect 14972 6500 14976 6556
rect 14976 6500 15032 6556
rect 15032 6500 15036 6556
rect 14972 6496 15036 6500
rect 20652 6556 20716 6560
rect 20652 6500 20656 6556
rect 20656 6500 20712 6556
rect 20712 6500 20716 6556
rect 20652 6496 20716 6500
rect 20732 6556 20796 6560
rect 20732 6500 20736 6556
rect 20736 6500 20792 6556
rect 20792 6500 20796 6556
rect 20732 6496 20796 6500
rect 20812 6556 20876 6560
rect 20812 6500 20816 6556
rect 20816 6500 20872 6556
rect 20872 6500 20876 6556
rect 20812 6496 20876 6500
rect 20892 6556 20956 6560
rect 20892 6500 20896 6556
rect 20896 6500 20952 6556
rect 20952 6500 20956 6556
rect 20892 6496 20956 6500
rect 20972 6556 21036 6560
rect 20972 6500 20976 6556
rect 20976 6500 21032 6556
rect 21032 6500 21036 6556
rect 20972 6496 21036 6500
rect 1912 6012 1976 6016
rect 1912 5956 1916 6012
rect 1916 5956 1972 6012
rect 1972 5956 1976 6012
rect 1912 5952 1976 5956
rect 1992 6012 2056 6016
rect 1992 5956 1996 6012
rect 1996 5956 2052 6012
rect 2052 5956 2056 6012
rect 1992 5952 2056 5956
rect 2072 6012 2136 6016
rect 2072 5956 2076 6012
rect 2076 5956 2132 6012
rect 2132 5956 2136 6012
rect 2072 5952 2136 5956
rect 2152 6012 2216 6016
rect 2152 5956 2156 6012
rect 2156 5956 2212 6012
rect 2212 5956 2216 6012
rect 2152 5952 2216 5956
rect 2232 6012 2296 6016
rect 2232 5956 2236 6012
rect 2236 5956 2292 6012
rect 2292 5956 2296 6012
rect 2232 5952 2296 5956
rect 7912 6012 7976 6016
rect 7912 5956 7916 6012
rect 7916 5956 7972 6012
rect 7972 5956 7976 6012
rect 7912 5952 7976 5956
rect 7992 6012 8056 6016
rect 7992 5956 7996 6012
rect 7996 5956 8052 6012
rect 8052 5956 8056 6012
rect 7992 5952 8056 5956
rect 8072 6012 8136 6016
rect 8072 5956 8076 6012
rect 8076 5956 8132 6012
rect 8132 5956 8136 6012
rect 8072 5952 8136 5956
rect 8152 6012 8216 6016
rect 8152 5956 8156 6012
rect 8156 5956 8212 6012
rect 8212 5956 8216 6012
rect 8152 5952 8216 5956
rect 8232 6012 8296 6016
rect 8232 5956 8236 6012
rect 8236 5956 8292 6012
rect 8292 5956 8296 6012
rect 8232 5952 8296 5956
rect 13912 6012 13976 6016
rect 13912 5956 13916 6012
rect 13916 5956 13972 6012
rect 13972 5956 13976 6012
rect 13912 5952 13976 5956
rect 13992 6012 14056 6016
rect 13992 5956 13996 6012
rect 13996 5956 14052 6012
rect 14052 5956 14056 6012
rect 13992 5952 14056 5956
rect 14072 6012 14136 6016
rect 14072 5956 14076 6012
rect 14076 5956 14132 6012
rect 14132 5956 14136 6012
rect 14072 5952 14136 5956
rect 14152 6012 14216 6016
rect 14152 5956 14156 6012
rect 14156 5956 14212 6012
rect 14212 5956 14216 6012
rect 14152 5952 14216 5956
rect 14232 6012 14296 6016
rect 14232 5956 14236 6012
rect 14236 5956 14292 6012
rect 14292 5956 14296 6012
rect 14232 5952 14296 5956
rect 19912 6012 19976 6016
rect 19912 5956 19916 6012
rect 19916 5956 19972 6012
rect 19972 5956 19976 6012
rect 19912 5952 19976 5956
rect 19992 6012 20056 6016
rect 19992 5956 19996 6012
rect 19996 5956 20052 6012
rect 20052 5956 20056 6012
rect 19992 5952 20056 5956
rect 20072 6012 20136 6016
rect 20072 5956 20076 6012
rect 20076 5956 20132 6012
rect 20132 5956 20136 6012
rect 20072 5952 20136 5956
rect 20152 6012 20216 6016
rect 20152 5956 20156 6012
rect 20156 5956 20212 6012
rect 20212 5956 20216 6012
rect 20152 5952 20216 5956
rect 20232 6012 20296 6016
rect 20232 5956 20236 6012
rect 20236 5956 20292 6012
rect 20292 5956 20296 6012
rect 20232 5952 20296 5956
rect 2652 5468 2716 5472
rect 2652 5412 2656 5468
rect 2656 5412 2712 5468
rect 2712 5412 2716 5468
rect 2652 5408 2716 5412
rect 2732 5468 2796 5472
rect 2732 5412 2736 5468
rect 2736 5412 2792 5468
rect 2792 5412 2796 5468
rect 2732 5408 2796 5412
rect 2812 5468 2876 5472
rect 2812 5412 2816 5468
rect 2816 5412 2872 5468
rect 2872 5412 2876 5468
rect 2812 5408 2876 5412
rect 2892 5468 2956 5472
rect 2892 5412 2896 5468
rect 2896 5412 2952 5468
rect 2952 5412 2956 5468
rect 2892 5408 2956 5412
rect 2972 5468 3036 5472
rect 2972 5412 2976 5468
rect 2976 5412 3032 5468
rect 3032 5412 3036 5468
rect 2972 5408 3036 5412
rect 8652 5468 8716 5472
rect 8652 5412 8656 5468
rect 8656 5412 8712 5468
rect 8712 5412 8716 5468
rect 8652 5408 8716 5412
rect 8732 5468 8796 5472
rect 8732 5412 8736 5468
rect 8736 5412 8792 5468
rect 8792 5412 8796 5468
rect 8732 5408 8796 5412
rect 8812 5468 8876 5472
rect 8812 5412 8816 5468
rect 8816 5412 8872 5468
rect 8872 5412 8876 5468
rect 8812 5408 8876 5412
rect 8892 5468 8956 5472
rect 8892 5412 8896 5468
rect 8896 5412 8952 5468
rect 8952 5412 8956 5468
rect 8892 5408 8956 5412
rect 8972 5468 9036 5472
rect 8972 5412 8976 5468
rect 8976 5412 9032 5468
rect 9032 5412 9036 5468
rect 8972 5408 9036 5412
rect 14652 5468 14716 5472
rect 14652 5412 14656 5468
rect 14656 5412 14712 5468
rect 14712 5412 14716 5468
rect 14652 5408 14716 5412
rect 14732 5468 14796 5472
rect 14732 5412 14736 5468
rect 14736 5412 14792 5468
rect 14792 5412 14796 5468
rect 14732 5408 14796 5412
rect 14812 5468 14876 5472
rect 14812 5412 14816 5468
rect 14816 5412 14872 5468
rect 14872 5412 14876 5468
rect 14812 5408 14876 5412
rect 14892 5468 14956 5472
rect 14892 5412 14896 5468
rect 14896 5412 14952 5468
rect 14952 5412 14956 5468
rect 14892 5408 14956 5412
rect 14972 5468 15036 5472
rect 14972 5412 14976 5468
rect 14976 5412 15032 5468
rect 15032 5412 15036 5468
rect 14972 5408 15036 5412
rect 20652 5468 20716 5472
rect 20652 5412 20656 5468
rect 20656 5412 20712 5468
rect 20712 5412 20716 5468
rect 20652 5408 20716 5412
rect 20732 5468 20796 5472
rect 20732 5412 20736 5468
rect 20736 5412 20792 5468
rect 20792 5412 20796 5468
rect 20732 5408 20796 5412
rect 20812 5468 20876 5472
rect 20812 5412 20816 5468
rect 20816 5412 20872 5468
rect 20872 5412 20876 5468
rect 20812 5408 20876 5412
rect 20892 5468 20956 5472
rect 20892 5412 20896 5468
rect 20896 5412 20952 5468
rect 20952 5412 20956 5468
rect 20892 5408 20956 5412
rect 20972 5468 21036 5472
rect 20972 5412 20976 5468
rect 20976 5412 21032 5468
rect 21032 5412 21036 5468
rect 20972 5408 21036 5412
rect 1912 4924 1976 4928
rect 1912 4868 1916 4924
rect 1916 4868 1972 4924
rect 1972 4868 1976 4924
rect 1912 4864 1976 4868
rect 1992 4924 2056 4928
rect 1992 4868 1996 4924
rect 1996 4868 2052 4924
rect 2052 4868 2056 4924
rect 1992 4864 2056 4868
rect 2072 4924 2136 4928
rect 2072 4868 2076 4924
rect 2076 4868 2132 4924
rect 2132 4868 2136 4924
rect 2072 4864 2136 4868
rect 2152 4924 2216 4928
rect 2152 4868 2156 4924
rect 2156 4868 2212 4924
rect 2212 4868 2216 4924
rect 2152 4864 2216 4868
rect 2232 4924 2296 4928
rect 2232 4868 2236 4924
rect 2236 4868 2292 4924
rect 2292 4868 2296 4924
rect 2232 4864 2296 4868
rect 7912 4924 7976 4928
rect 7912 4868 7916 4924
rect 7916 4868 7972 4924
rect 7972 4868 7976 4924
rect 7912 4864 7976 4868
rect 7992 4924 8056 4928
rect 7992 4868 7996 4924
rect 7996 4868 8052 4924
rect 8052 4868 8056 4924
rect 7992 4864 8056 4868
rect 8072 4924 8136 4928
rect 8072 4868 8076 4924
rect 8076 4868 8132 4924
rect 8132 4868 8136 4924
rect 8072 4864 8136 4868
rect 8152 4924 8216 4928
rect 8152 4868 8156 4924
rect 8156 4868 8212 4924
rect 8212 4868 8216 4924
rect 8152 4864 8216 4868
rect 8232 4924 8296 4928
rect 8232 4868 8236 4924
rect 8236 4868 8292 4924
rect 8292 4868 8296 4924
rect 8232 4864 8296 4868
rect 13912 4924 13976 4928
rect 13912 4868 13916 4924
rect 13916 4868 13972 4924
rect 13972 4868 13976 4924
rect 13912 4864 13976 4868
rect 13992 4924 14056 4928
rect 13992 4868 13996 4924
rect 13996 4868 14052 4924
rect 14052 4868 14056 4924
rect 13992 4864 14056 4868
rect 14072 4924 14136 4928
rect 14072 4868 14076 4924
rect 14076 4868 14132 4924
rect 14132 4868 14136 4924
rect 14072 4864 14136 4868
rect 14152 4924 14216 4928
rect 14152 4868 14156 4924
rect 14156 4868 14212 4924
rect 14212 4868 14216 4924
rect 14152 4864 14216 4868
rect 14232 4924 14296 4928
rect 14232 4868 14236 4924
rect 14236 4868 14292 4924
rect 14292 4868 14296 4924
rect 14232 4864 14296 4868
rect 19912 4924 19976 4928
rect 19912 4868 19916 4924
rect 19916 4868 19972 4924
rect 19972 4868 19976 4924
rect 19912 4864 19976 4868
rect 19992 4924 20056 4928
rect 19992 4868 19996 4924
rect 19996 4868 20052 4924
rect 20052 4868 20056 4924
rect 19992 4864 20056 4868
rect 20072 4924 20136 4928
rect 20072 4868 20076 4924
rect 20076 4868 20132 4924
rect 20132 4868 20136 4924
rect 20072 4864 20136 4868
rect 20152 4924 20216 4928
rect 20152 4868 20156 4924
rect 20156 4868 20212 4924
rect 20212 4868 20216 4924
rect 20152 4864 20216 4868
rect 20232 4924 20296 4928
rect 20232 4868 20236 4924
rect 20236 4868 20292 4924
rect 20292 4868 20296 4924
rect 20232 4864 20296 4868
rect 2652 4380 2716 4384
rect 2652 4324 2656 4380
rect 2656 4324 2712 4380
rect 2712 4324 2716 4380
rect 2652 4320 2716 4324
rect 2732 4380 2796 4384
rect 2732 4324 2736 4380
rect 2736 4324 2792 4380
rect 2792 4324 2796 4380
rect 2732 4320 2796 4324
rect 2812 4380 2876 4384
rect 2812 4324 2816 4380
rect 2816 4324 2872 4380
rect 2872 4324 2876 4380
rect 2812 4320 2876 4324
rect 2892 4380 2956 4384
rect 2892 4324 2896 4380
rect 2896 4324 2952 4380
rect 2952 4324 2956 4380
rect 2892 4320 2956 4324
rect 2972 4380 3036 4384
rect 2972 4324 2976 4380
rect 2976 4324 3032 4380
rect 3032 4324 3036 4380
rect 2972 4320 3036 4324
rect 8652 4380 8716 4384
rect 8652 4324 8656 4380
rect 8656 4324 8712 4380
rect 8712 4324 8716 4380
rect 8652 4320 8716 4324
rect 8732 4380 8796 4384
rect 8732 4324 8736 4380
rect 8736 4324 8792 4380
rect 8792 4324 8796 4380
rect 8732 4320 8796 4324
rect 8812 4380 8876 4384
rect 8812 4324 8816 4380
rect 8816 4324 8872 4380
rect 8872 4324 8876 4380
rect 8812 4320 8876 4324
rect 8892 4380 8956 4384
rect 8892 4324 8896 4380
rect 8896 4324 8952 4380
rect 8952 4324 8956 4380
rect 8892 4320 8956 4324
rect 8972 4380 9036 4384
rect 8972 4324 8976 4380
rect 8976 4324 9032 4380
rect 9032 4324 9036 4380
rect 8972 4320 9036 4324
rect 14652 4380 14716 4384
rect 14652 4324 14656 4380
rect 14656 4324 14712 4380
rect 14712 4324 14716 4380
rect 14652 4320 14716 4324
rect 14732 4380 14796 4384
rect 14732 4324 14736 4380
rect 14736 4324 14792 4380
rect 14792 4324 14796 4380
rect 14732 4320 14796 4324
rect 14812 4380 14876 4384
rect 14812 4324 14816 4380
rect 14816 4324 14872 4380
rect 14872 4324 14876 4380
rect 14812 4320 14876 4324
rect 14892 4380 14956 4384
rect 14892 4324 14896 4380
rect 14896 4324 14952 4380
rect 14952 4324 14956 4380
rect 14892 4320 14956 4324
rect 14972 4380 15036 4384
rect 14972 4324 14976 4380
rect 14976 4324 15032 4380
rect 15032 4324 15036 4380
rect 14972 4320 15036 4324
rect 20652 4380 20716 4384
rect 20652 4324 20656 4380
rect 20656 4324 20712 4380
rect 20712 4324 20716 4380
rect 20652 4320 20716 4324
rect 20732 4380 20796 4384
rect 20732 4324 20736 4380
rect 20736 4324 20792 4380
rect 20792 4324 20796 4380
rect 20732 4320 20796 4324
rect 20812 4380 20876 4384
rect 20812 4324 20816 4380
rect 20816 4324 20872 4380
rect 20872 4324 20876 4380
rect 20812 4320 20876 4324
rect 20892 4380 20956 4384
rect 20892 4324 20896 4380
rect 20896 4324 20952 4380
rect 20952 4324 20956 4380
rect 20892 4320 20956 4324
rect 20972 4380 21036 4384
rect 20972 4324 20976 4380
rect 20976 4324 21032 4380
rect 21032 4324 21036 4380
rect 20972 4320 21036 4324
rect 1912 3836 1976 3840
rect 1912 3780 1916 3836
rect 1916 3780 1972 3836
rect 1972 3780 1976 3836
rect 1912 3776 1976 3780
rect 1992 3836 2056 3840
rect 1992 3780 1996 3836
rect 1996 3780 2052 3836
rect 2052 3780 2056 3836
rect 1992 3776 2056 3780
rect 2072 3836 2136 3840
rect 2072 3780 2076 3836
rect 2076 3780 2132 3836
rect 2132 3780 2136 3836
rect 2072 3776 2136 3780
rect 2152 3836 2216 3840
rect 2152 3780 2156 3836
rect 2156 3780 2212 3836
rect 2212 3780 2216 3836
rect 2152 3776 2216 3780
rect 2232 3836 2296 3840
rect 2232 3780 2236 3836
rect 2236 3780 2292 3836
rect 2292 3780 2296 3836
rect 2232 3776 2296 3780
rect 7912 3836 7976 3840
rect 7912 3780 7916 3836
rect 7916 3780 7972 3836
rect 7972 3780 7976 3836
rect 7912 3776 7976 3780
rect 7992 3836 8056 3840
rect 7992 3780 7996 3836
rect 7996 3780 8052 3836
rect 8052 3780 8056 3836
rect 7992 3776 8056 3780
rect 8072 3836 8136 3840
rect 8072 3780 8076 3836
rect 8076 3780 8132 3836
rect 8132 3780 8136 3836
rect 8072 3776 8136 3780
rect 8152 3836 8216 3840
rect 8152 3780 8156 3836
rect 8156 3780 8212 3836
rect 8212 3780 8216 3836
rect 8152 3776 8216 3780
rect 8232 3836 8296 3840
rect 8232 3780 8236 3836
rect 8236 3780 8292 3836
rect 8292 3780 8296 3836
rect 8232 3776 8296 3780
rect 13912 3836 13976 3840
rect 13912 3780 13916 3836
rect 13916 3780 13972 3836
rect 13972 3780 13976 3836
rect 13912 3776 13976 3780
rect 13992 3836 14056 3840
rect 13992 3780 13996 3836
rect 13996 3780 14052 3836
rect 14052 3780 14056 3836
rect 13992 3776 14056 3780
rect 14072 3836 14136 3840
rect 14072 3780 14076 3836
rect 14076 3780 14132 3836
rect 14132 3780 14136 3836
rect 14072 3776 14136 3780
rect 14152 3836 14216 3840
rect 14152 3780 14156 3836
rect 14156 3780 14212 3836
rect 14212 3780 14216 3836
rect 14152 3776 14216 3780
rect 14232 3836 14296 3840
rect 14232 3780 14236 3836
rect 14236 3780 14292 3836
rect 14292 3780 14296 3836
rect 14232 3776 14296 3780
rect 19912 3836 19976 3840
rect 19912 3780 19916 3836
rect 19916 3780 19972 3836
rect 19972 3780 19976 3836
rect 19912 3776 19976 3780
rect 19992 3836 20056 3840
rect 19992 3780 19996 3836
rect 19996 3780 20052 3836
rect 20052 3780 20056 3836
rect 19992 3776 20056 3780
rect 20072 3836 20136 3840
rect 20072 3780 20076 3836
rect 20076 3780 20132 3836
rect 20132 3780 20136 3836
rect 20072 3776 20136 3780
rect 20152 3836 20216 3840
rect 20152 3780 20156 3836
rect 20156 3780 20212 3836
rect 20212 3780 20216 3836
rect 20152 3776 20216 3780
rect 20232 3836 20296 3840
rect 20232 3780 20236 3836
rect 20236 3780 20292 3836
rect 20292 3780 20296 3836
rect 20232 3776 20296 3780
rect 2652 3292 2716 3296
rect 2652 3236 2656 3292
rect 2656 3236 2712 3292
rect 2712 3236 2716 3292
rect 2652 3232 2716 3236
rect 2732 3292 2796 3296
rect 2732 3236 2736 3292
rect 2736 3236 2792 3292
rect 2792 3236 2796 3292
rect 2732 3232 2796 3236
rect 2812 3292 2876 3296
rect 2812 3236 2816 3292
rect 2816 3236 2872 3292
rect 2872 3236 2876 3292
rect 2812 3232 2876 3236
rect 2892 3292 2956 3296
rect 2892 3236 2896 3292
rect 2896 3236 2952 3292
rect 2952 3236 2956 3292
rect 2892 3232 2956 3236
rect 2972 3292 3036 3296
rect 2972 3236 2976 3292
rect 2976 3236 3032 3292
rect 3032 3236 3036 3292
rect 2972 3232 3036 3236
rect 8652 3292 8716 3296
rect 8652 3236 8656 3292
rect 8656 3236 8712 3292
rect 8712 3236 8716 3292
rect 8652 3232 8716 3236
rect 8732 3292 8796 3296
rect 8732 3236 8736 3292
rect 8736 3236 8792 3292
rect 8792 3236 8796 3292
rect 8732 3232 8796 3236
rect 8812 3292 8876 3296
rect 8812 3236 8816 3292
rect 8816 3236 8872 3292
rect 8872 3236 8876 3292
rect 8812 3232 8876 3236
rect 8892 3292 8956 3296
rect 8892 3236 8896 3292
rect 8896 3236 8952 3292
rect 8952 3236 8956 3292
rect 8892 3232 8956 3236
rect 8972 3292 9036 3296
rect 8972 3236 8976 3292
rect 8976 3236 9032 3292
rect 9032 3236 9036 3292
rect 8972 3232 9036 3236
rect 14652 3292 14716 3296
rect 14652 3236 14656 3292
rect 14656 3236 14712 3292
rect 14712 3236 14716 3292
rect 14652 3232 14716 3236
rect 14732 3292 14796 3296
rect 14732 3236 14736 3292
rect 14736 3236 14792 3292
rect 14792 3236 14796 3292
rect 14732 3232 14796 3236
rect 14812 3292 14876 3296
rect 14812 3236 14816 3292
rect 14816 3236 14872 3292
rect 14872 3236 14876 3292
rect 14812 3232 14876 3236
rect 14892 3292 14956 3296
rect 14892 3236 14896 3292
rect 14896 3236 14952 3292
rect 14952 3236 14956 3292
rect 14892 3232 14956 3236
rect 14972 3292 15036 3296
rect 14972 3236 14976 3292
rect 14976 3236 15032 3292
rect 15032 3236 15036 3292
rect 14972 3232 15036 3236
rect 20652 3292 20716 3296
rect 20652 3236 20656 3292
rect 20656 3236 20712 3292
rect 20712 3236 20716 3292
rect 20652 3232 20716 3236
rect 20732 3292 20796 3296
rect 20732 3236 20736 3292
rect 20736 3236 20792 3292
rect 20792 3236 20796 3292
rect 20732 3232 20796 3236
rect 20812 3292 20876 3296
rect 20812 3236 20816 3292
rect 20816 3236 20872 3292
rect 20872 3236 20876 3292
rect 20812 3232 20876 3236
rect 20892 3292 20956 3296
rect 20892 3236 20896 3292
rect 20896 3236 20952 3292
rect 20952 3236 20956 3292
rect 20892 3232 20956 3236
rect 20972 3292 21036 3296
rect 20972 3236 20976 3292
rect 20976 3236 21032 3292
rect 21032 3236 21036 3292
rect 20972 3232 21036 3236
rect 1912 2748 1976 2752
rect 1912 2692 1916 2748
rect 1916 2692 1972 2748
rect 1972 2692 1976 2748
rect 1912 2688 1976 2692
rect 1992 2748 2056 2752
rect 1992 2692 1996 2748
rect 1996 2692 2052 2748
rect 2052 2692 2056 2748
rect 1992 2688 2056 2692
rect 2072 2748 2136 2752
rect 2072 2692 2076 2748
rect 2076 2692 2132 2748
rect 2132 2692 2136 2748
rect 2072 2688 2136 2692
rect 2152 2748 2216 2752
rect 2152 2692 2156 2748
rect 2156 2692 2212 2748
rect 2212 2692 2216 2748
rect 2152 2688 2216 2692
rect 2232 2748 2296 2752
rect 2232 2692 2236 2748
rect 2236 2692 2292 2748
rect 2292 2692 2296 2748
rect 2232 2688 2296 2692
rect 7912 2748 7976 2752
rect 7912 2692 7916 2748
rect 7916 2692 7972 2748
rect 7972 2692 7976 2748
rect 7912 2688 7976 2692
rect 7992 2748 8056 2752
rect 7992 2692 7996 2748
rect 7996 2692 8052 2748
rect 8052 2692 8056 2748
rect 7992 2688 8056 2692
rect 8072 2748 8136 2752
rect 8072 2692 8076 2748
rect 8076 2692 8132 2748
rect 8132 2692 8136 2748
rect 8072 2688 8136 2692
rect 8152 2748 8216 2752
rect 8152 2692 8156 2748
rect 8156 2692 8212 2748
rect 8212 2692 8216 2748
rect 8152 2688 8216 2692
rect 8232 2748 8296 2752
rect 8232 2692 8236 2748
rect 8236 2692 8292 2748
rect 8292 2692 8296 2748
rect 8232 2688 8296 2692
rect 13912 2748 13976 2752
rect 13912 2692 13916 2748
rect 13916 2692 13972 2748
rect 13972 2692 13976 2748
rect 13912 2688 13976 2692
rect 13992 2748 14056 2752
rect 13992 2692 13996 2748
rect 13996 2692 14052 2748
rect 14052 2692 14056 2748
rect 13992 2688 14056 2692
rect 14072 2748 14136 2752
rect 14072 2692 14076 2748
rect 14076 2692 14132 2748
rect 14132 2692 14136 2748
rect 14072 2688 14136 2692
rect 14152 2748 14216 2752
rect 14152 2692 14156 2748
rect 14156 2692 14212 2748
rect 14212 2692 14216 2748
rect 14152 2688 14216 2692
rect 14232 2748 14296 2752
rect 14232 2692 14236 2748
rect 14236 2692 14292 2748
rect 14292 2692 14296 2748
rect 14232 2688 14296 2692
rect 19912 2748 19976 2752
rect 19912 2692 19916 2748
rect 19916 2692 19972 2748
rect 19972 2692 19976 2748
rect 19912 2688 19976 2692
rect 19992 2748 20056 2752
rect 19992 2692 19996 2748
rect 19996 2692 20052 2748
rect 20052 2692 20056 2748
rect 19992 2688 20056 2692
rect 20072 2748 20136 2752
rect 20072 2692 20076 2748
rect 20076 2692 20132 2748
rect 20132 2692 20136 2748
rect 20072 2688 20136 2692
rect 20152 2748 20216 2752
rect 20152 2692 20156 2748
rect 20156 2692 20212 2748
rect 20212 2692 20216 2748
rect 20152 2688 20216 2692
rect 20232 2748 20296 2752
rect 20232 2692 20236 2748
rect 20236 2692 20292 2748
rect 20292 2692 20296 2748
rect 20232 2688 20296 2692
rect 2652 2204 2716 2208
rect 2652 2148 2656 2204
rect 2656 2148 2712 2204
rect 2712 2148 2716 2204
rect 2652 2144 2716 2148
rect 2732 2204 2796 2208
rect 2732 2148 2736 2204
rect 2736 2148 2792 2204
rect 2792 2148 2796 2204
rect 2732 2144 2796 2148
rect 2812 2204 2876 2208
rect 2812 2148 2816 2204
rect 2816 2148 2872 2204
rect 2872 2148 2876 2204
rect 2812 2144 2876 2148
rect 2892 2204 2956 2208
rect 2892 2148 2896 2204
rect 2896 2148 2952 2204
rect 2952 2148 2956 2204
rect 2892 2144 2956 2148
rect 2972 2204 3036 2208
rect 2972 2148 2976 2204
rect 2976 2148 3032 2204
rect 3032 2148 3036 2204
rect 2972 2144 3036 2148
rect 8652 2204 8716 2208
rect 8652 2148 8656 2204
rect 8656 2148 8712 2204
rect 8712 2148 8716 2204
rect 8652 2144 8716 2148
rect 8732 2204 8796 2208
rect 8732 2148 8736 2204
rect 8736 2148 8792 2204
rect 8792 2148 8796 2204
rect 8732 2144 8796 2148
rect 8812 2204 8876 2208
rect 8812 2148 8816 2204
rect 8816 2148 8872 2204
rect 8872 2148 8876 2204
rect 8812 2144 8876 2148
rect 8892 2204 8956 2208
rect 8892 2148 8896 2204
rect 8896 2148 8952 2204
rect 8952 2148 8956 2204
rect 8892 2144 8956 2148
rect 8972 2204 9036 2208
rect 8972 2148 8976 2204
rect 8976 2148 9032 2204
rect 9032 2148 9036 2204
rect 8972 2144 9036 2148
rect 14652 2204 14716 2208
rect 14652 2148 14656 2204
rect 14656 2148 14712 2204
rect 14712 2148 14716 2204
rect 14652 2144 14716 2148
rect 14732 2204 14796 2208
rect 14732 2148 14736 2204
rect 14736 2148 14792 2204
rect 14792 2148 14796 2204
rect 14732 2144 14796 2148
rect 14812 2204 14876 2208
rect 14812 2148 14816 2204
rect 14816 2148 14872 2204
rect 14872 2148 14876 2204
rect 14812 2144 14876 2148
rect 14892 2204 14956 2208
rect 14892 2148 14896 2204
rect 14896 2148 14952 2204
rect 14952 2148 14956 2204
rect 14892 2144 14956 2148
rect 14972 2204 15036 2208
rect 14972 2148 14976 2204
rect 14976 2148 15032 2204
rect 15032 2148 15036 2204
rect 14972 2144 15036 2148
rect 20652 2204 20716 2208
rect 20652 2148 20656 2204
rect 20656 2148 20712 2204
rect 20712 2148 20716 2204
rect 20652 2144 20716 2148
rect 20732 2204 20796 2208
rect 20732 2148 20736 2204
rect 20736 2148 20792 2204
rect 20792 2148 20796 2204
rect 20732 2144 20796 2148
rect 20812 2204 20876 2208
rect 20812 2148 20816 2204
rect 20816 2148 20872 2204
rect 20872 2148 20876 2204
rect 20812 2144 20876 2148
rect 20892 2204 20956 2208
rect 20892 2148 20896 2204
rect 20896 2148 20952 2204
rect 20952 2148 20956 2204
rect 20892 2144 20956 2148
rect 20972 2204 21036 2208
rect 20972 2148 20976 2204
rect 20976 2148 21032 2204
rect 21032 2148 21036 2204
rect 20972 2144 21036 2148
<< metal4 >>
rect -1076 26618 -756 26660
rect -1076 26382 -1034 26618
rect -798 26382 -756 26618
rect -1076 22034 -756 26382
rect -1076 21798 -1034 22034
rect -798 21798 -756 22034
rect -1076 16034 -756 21798
rect -1076 15798 -1034 16034
rect -798 15798 -756 16034
rect -1076 10034 -756 15798
rect -1076 9798 -1034 10034
rect -798 9798 -756 10034
rect -1076 4034 -756 9798
rect -1076 3798 -1034 4034
rect -798 3798 -756 4034
rect -1076 274 -756 3798
rect -416 25958 -96 26000
rect -416 25722 -374 25958
rect -138 25722 -96 25958
rect -416 21294 -96 25722
rect -416 21058 -374 21294
rect -138 21058 -96 21294
rect -416 15294 -96 21058
rect -416 15058 -374 15294
rect -138 15058 -96 15294
rect -416 9294 -96 15058
rect -416 9058 -374 9294
rect -138 9058 -96 9294
rect -416 3294 -96 9058
rect -416 3058 -374 3294
rect -138 3058 -96 3294
rect -416 934 -96 3058
rect -416 698 -374 934
rect -138 698 -96 934
rect -416 656 -96 698
rect 1904 25958 2304 26660
rect 1904 25722 1986 25958
rect 2222 25722 2304 25958
rect 1904 24512 2304 25722
rect 1904 24448 1912 24512
rect 1976 24448 1992 24512
rect 2056 24448 2072 24512
rect 2136 24448 2152 24512
rect 2216 24448 2232 24512
rect 2296 24448 2304 24512
rect 1904 23424 2304 24448
rect 1904 23360 1912 23424
rect 1976 23360 1992 23424
rect 2056 23360 2072 23424
rect 2136 23360 2152 23424
rect 2216 23360 2232 23424
rect 2296 23360 2304 23424
rect 1904 22336 2304 23360
rect 1904 22272 1912 22336
rect 1976 22272 1992 22336
rect 2056 22272 2072 22336
rect 2136 22272 2152 22336
rect 2216 22272 2232 22336
rect 2296 22272 2304 22336
rect 1904 21294 2304 22272
rect 1904 21248 1986 21294
rect 2222 21248 2304 21294
rect 1904 21184 1912 21248
rect 1976 21184 1986 21248
rect 2222 21184 2232 21248
rect 2296 21184 2304 21248
rect 1904 21058 1986 21184
rect 2222 21058 2304 21184
rect 1904 20160 2304 21058
rect 1904 20096 1912 20160
rect 1976 20096 1992 20160
rect 2056 20096 2072 20160
rect 2136 20096 2152 20160
rect 2216 20096 2232 20160
rect 2296 20096 2304 20160
rect 1904 19072 2304 20096
rect 1904 19008 1912 19072
rect 1976 19008 1992 19072
rect 2056 19008 2072 19072
rect 2136 19008 2152 19072
rect 2216 19008 2232 19072
rect 2296 19008 2304 19072
rect 1904 17984 2304 19008
rect 1904 17920 1912 17984
rect 1976 17920 1992 17984
rect 2056 17920 2072 17984
rect 2136 17920 2152 17984
rect 2216 17920 2232 17984
rect 2296 17920 2304 17984
rect 1904 16896 2304 17920
rect 1904 16832 1912 16896
rect 1976 16832 1992 16896
rect 2056 16832 2072 16896
rect 2136 16832 2152 16896
rect 2216 16832 2232 16896
rect 2296 16832 2304 16896
rect 1904 15808 2304 16832
rect 1904 15744 1912 15808
rect 1976 15744 1992 15808
rect 2056 15744 2072 15808
rect 2136 15744 2152 15808
rect 2216 15744 2232 15808
rect 2296 15744 2304 15808
rect 1904 15294 2304 15744
rect 1904 15058 1986 15294
rect 2222 15058 2304 15294
rect 1904 14720 2304 15058
rect 1904 14656 1912 14720
rect 1976 14656 1992 14720
rect 2056 14656 2072 14720
rect 2136 14656 2152 14720
rect 2216 14656 2232 14720
rect 2296 14656 2304 14720
rect 1904 13632 2304 14656
rect 1904 13568 1912 13632
rect 1976 13568 1992 13632
rect 2056 13568 2072 13632
rect 2136 13568 2152 13632
rect 2216 13568 2232 13632
rect 2296 13568 2304 13632
rect 1904 12544 2304 13568
rect 1904 12480 1912 12544
rect 1976 12480 1992 12544
rect 2056 12480 2072 12544
rect 2136 12480 2152 12544
rect 2216 12480 2232 12544
rect 2296 12480 2304 12544
rect 1904 11456 2304 12480
rect 1904 11392 1912 11456
rect 1976 11392 1992 11456
rect 2056 11392 2072 11456
rect 2136 11392 2152 11456
rect 2216 11392 2232 11456
rect 2296 11392 2304 11456
rect 1904 10368 2304 11392
rect 1904 10304 1912 10368
rect 1976 10304 1992 10368
rect 2056 10304 2072 10368
rect 2136 10304 2152 10368
rect 2216 10304 2232 10368
rect 2296 10304 2304 10368
rect 1904 9294 2304 10304
rect 1904 9280 1986 9294
rect 2222 9280 2304 9294
rect 1904 9216 1912 9280
rect 1976 9216 1986 9280
rect 2222 9216 2232 9280
rect 2296 9216 2304 9280
rect 1904 9058 1986 9216
rect 2222 9058 2304 9216
rect 1904 8192 2304 9058
rect 1904 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2304 8192
rect 1904 7104 2304 8128
rect 1904 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2304 7104
rect 1904 6016 2304 7040
rect 1904 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2304 6016
rect 1904 4928 2304 5952
rect 1904 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2304 4928
rect 1904 3840 2304 4864
rect 1904 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2304 3840
rect 1904 3294 2304 3776
rect 1904 3058 1986 3294
rect 2222 3058 2304 3294
rect 1904 2752 2304 3058
rect 1904 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2304 2752
rect 1904 934 2304 2688
rect 1904 698 1986 934
rect 2222 698 2304 934
rect -1076 38 -1034 274
rect -798 38 -756 274
rect -1076 -4 -756 38
rect 1904 -4 2304 698
rect 2644 26618 3044 26660
rect 2644 26382 2726 26618
rect 2962 26382 3044 26618
rect 2644 23968 3044 26382
rect 2644 23904 2652 23968
rect 2716 23904 2732 23968
rect 2796 23904 2812 23968
rect 2876 23904 2892 23968
rect 2956 23904 2972 23968
rect 3036 23904 3044 23968
rect 2644 22880 3044 23904
rect 2644 22816 2652 22880
rect 2716 22816 2732 22880
rect 2796 22816 2812 22880
rect 2876 22816 2892 22880
rect 2956 22816 2972 22880
rect 3036 22816 3044 22880
rect 2644 22034 3044 22816
rect 2644 21798 2726 22034
rect 2962 21798 3044 22034
rect 2644 21792 3044 21798
rect 2644 21728 2652 21792
rect 2716 21728 2732 21792
rect 2796 21728 2812 21792
rect 2876 21728 2892 21792
rect 2956 21728 2972 21792
rect 3036 21728 3044 21792
rect 2644 20704 3044 21728
rect 2644 20640 2652 20704
rect 2716 20640 2732 20704
rect 2796 20640 2812 20704
rect 2876 20640 2892 20704
rect 2956 20640 2972 20704
rect 3036 20640 3044 20704
rect 2644 19616 3044 20640
rect 2644 19552 2652 19616
rect 2716 19552 2732 19616
rect 2796 19552 2812 19616
rect 2876 19552 2892 19616
rect 2956 19552 2972 19616
rect 3036 19552 3044 19616
rect 2644 18528 3044 19552
rect 2644 18464 2652 18528
rect 2716 18464 2732 18528
rect 2796 18464 2812 18528
rect 2876 18464 2892 18528
rect 2956 18464 2972 18528
rect 3036 18464 3044 18528
rect 2644 17440 3044 18464
rect 2644 17376 2652 17440
rect 2716 17376 2732 17440
rect 2796 17376 2812 17440
rect 2876 17376 2892 17440
rect 2956 17376 2972 17440
rect 3036 17376 3044 17440
rect 2644 16352 3044 17376
rect 2644 16288 2652 16352
rect 2716 16288 2732 16352
rect 2796 16288 2812 16352
rect 2876 16288 2892 16352
rect 2956 16288 2972 16352
rect 3036 16288 3044 16352
rect 2644 16034 3044 16288
rect 2644 15798 2726 16034
rect 2962 15798 3044 16034
rect 2644 15264 3044 15798
rect 2644 15200 2652 15264
rect 2716 15200 2732 15264
rect 2796 15200 2812 15264
rect 2876 15200 2892 15264
rect 2956 15200 2972 15264
rect 3036 15200 3044 15264
rect 2644 14176 3044 15200
rect 2644 14112 2652 14176
rect 2716 14112 2732 14176
rect 2796 14112 2812 14176
rect 2876 14112 2892 14176
rect 2956 14112 2972 14176
rect 3036 14112 3044 14176
rect 2644 13088 3044 14112
rect 2644 13024 2652 13088
rect 2716 13024 2732 13088
rect 2796 13024 2812 13088
rect 2876 13024 2892 13088
rect 2956 13024 2972 13088
rect 3036 13024 3044 13088
rect 2644 12000 3044 13024
rect 2644 11936 2652 12000
rect 2716 11936 2732 12000
rect 2796 11936 2812 12000
rect 2876 11936 2892 12000
rect 2956 11936 2972 12000
rect 3036 11936 3044 12000
rect 2644 10912 3044 11936
rect 2644 10848 2652 10912
rect 2716 10848 2732 10912
rect 2796 10848 2812 10912
rect 2876 10848 2892 10912
rect 2956 10848 2972 10912
rect 3036 10848 3044 10912
rect 2644 10034 3044 10848
rect 2644 9824 2726 10034
rect 2962 9824 3044 10034
rect 2644 9760 2652 9824
rect 2716 9798 2726 9824
rect 2962 9798 2972 9824
rect 2716 9760 2732 9798
rect 2796 9760 2812 9798
rect 2876 9760 2892 9798
rect 2956 9760 2972 9798
rect 3036 9760 3044 9824
rect 2644 8736 3044 9760
rect 2644 8672 2652 8736
rect 2716 8672 2732 8736
rect 2796 8672 2812 8736
rect 2876 8672 2892 8736
rect 2956 8672 2972 8736
rect 3036 8672 3044 8736
rect 2644 7648 3044 8672
rect 2644 7584 2652 7648
rect 2716 7584 2732 7648
rect 2796 7584 2812 7648
rect 2876 7584 2892 7648
rect 2956 7584 2972 7648
rect 3036 7584 3044 7648
rect 2644 6560 3044 7584
rect 2644 6496 2652 6560
rect 2716 6496 2732 6560
rect 2796 6496 2812 6560
rect 2876 6496 2892 6560
rect 2956 6496 2972 6560
rect 3036 6496 3044 6560
rect 2644 5472 3044 6496
rect 2644 5408 2652 5472
rect 2716 5408 2732 5472
rect 2796 5408 2812 5472
rect 2876 5408 2892 5472
rect 2956 5408 2972 5472
rect 3036 5408 3044 5472
rect 2644 4384 3044 5408
rect 2644 4320 2652 4384
rect 2716 4320 2732 4384
rect 2796 4320 2812 4384
rect 2876 4320 2892 4384
rect 2956 4320 2972 4384
rect 3036 4320 3044 4384
rect 2644 4034 3044 4320
rect 2644 3798 2726 4034
rect 2962 3798 3044 4034
rect 2644 3296 3044 3798
rect 2644 3232 2652 3296
rect 2716 3232 2732 3296
rect 2796 3232 2812 3296
rect 2876 3232 2892 3296
rect 2956 3232 2972 3296
rect 3036 3232 3044 3296
rect 2644 2208 3044 3232
rect 2644 2144 2652 2208
rect 2716 2144 2732 2208
rect 2796 2144 2812 2208
rect 2876 2144 2892 2208
rect 2956 2144 2972 2208
rect 3036 2144 3044 2208
rect 2644 274 3044 2144
rect 2644 38 2726 274
rect 2962 38 3044 274
rect 2644 -4 3044 38
rect 7904 25958 8304 26660
rect 7904 25722 7986 25958
rect 8222 25722 8304 25958
rect 7904 24512 8304 25722
rect 7904 24448 7912 24512
rect 7976 24448 7992 24512
rect 8056 24448 8072 24512
rect 8136 24448 8152 24512
rect 8216 24448 8232 24512
rect 8296 24448 8304 24512
rect 7904 23424 8304 24448
rect 7904 23360 7912 23424
rect 7976 23360 7992 23424
rect 8056 23360 8072 23424
rect 8136 23360 8152 23424
rect 8216 23360 8232 23424
rect 8296 23360 8304 23424
rect 7904 22336 8304 23360
rect 7904 22272 7912 22336
rect 7976 22272 7992 22336
rect 8056 22272 8072 22336
rect 8136 22272 8152 22336
rect 8216 22272 8232 22336
rect 8296 22272 8304 22336
rect 7904 21294 8304 22272
rect 7904 21248 7986 21294
rect 8222 21248 8304 21294
rect 7904 21184 7912 21248
rect 7976 21184 7986 21248
rect 8222 21184 8232 21248
rect 8296 21184 8304 21248
rect 7904 21058 7986 21184
rect 8222 21058 8304 21184
rect 7904 20160 8304 21058
rect 7904 20096 7912 20160
rect 7976 20096 7992 20160
rect 8056 20096 8072 20160
rect 8136 20096 8152 20160
rect 8216 20096 8232 20160
rect 8296 20096 8304 20160
rect 7904 19072 8304 20096
rect 7904 19008 7912 19072
rect 7976 19008 7992 19072
rect 8056 19008 8072 19072
rect 8136 19008 8152 19072
rect 8216 19008 8232 19072
rect 8296 19008 8304 19072
rect 7904 17984 8304 19008
rect 7904 17920 7912 17984
rect 7976 17920 7992 17984
rect 8056 17920 8072 17984
rect 8136 17920 8152 17984
rect 8216 17920 8232 17984
rect 8296 17920 8304 17984
rect 7904 16896 8304 17920
rect 7904 16832 7912 16896
rect 7976 16832 7992 16896
rect 8056 16832 8072 16896
rect 8136 16832 8152 16896
rect 8216 16832 8232 16896
rect 8296 16832 8304 16896
rect 7904 15808 8304 16832
rect 7904 15744 7912 15808
rect 7976 15744 7992 15808
rect 8056 15744 8072 15808
rect 8136 15744 8152 15808
rect 8216 15744 8232 15808
rect 8296 15744 8304 15808
rect 7904 15294 8304 15744
rect 7904 15058 7986 15294
rect 8222 15058 8304 15294
rect 7904 14720 8304 15058
rect 7904 14656 7912 14720
rect 7976 14656 7992 14720
rect 8056 14656 8072 14720
rect 8136 14656 8152 14720
rect 8216 14656 8232 14720
rect 8296 14656 8304 14720
rect 7904 13632 8304 14656
rect 7904 13568 7912 13632
rect 7976 13568 7992 13632
rect 8056 13568 8072 13632
rect 8136 13568 8152 13632
rect 8216 13568 8232 13632
rect 8296 13568 8304 13632
rect 7904 12544 8304 13568
rect 7904 12480 7912 12544
rect 7976 12480 7992 12544
rect 8056 12480 8072 12544
rect 8136 12480 8152 12544
rect 8216 12480 8232 12544
rect 8296 12480 8304 12544
rect 7904 11456 8304 12480
rect 7904 11392 7912 11456
rect 7976 11392 7992 11456
rect 8056 11392 8072 11456
rect 8136 11392 8152 11456
rect 8216 11392 8232 11456
rect 8296 11392 8304 11456
rect 7904 10368 8304 11392
rect 7904 10304 7912 10368
rect 7976 10304 7992 10368
rect 8056 10304 8072 10368
rect 8136 10304 8152 10368
rect 8216 10304 8232 10368
rect 8296 10304 8304 10368
rect 7904 9294 8304 10304
rect 7904 9280 7986 9294
rect 8222 9280 8304 9294
rect 7904 9216 7912 9280
rect 7976 9216 7986 9280
rect 8222 9216 8232 9280
rect 8296 9216 8304 9280
rect 7904 9058 7986 9216
rect 8222 9058 8304 9216
rect 7904 8192 8304 9058
rect 7904 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8072 8192
rect 8136 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8304 8192
rect 7904 7104 8304 8128
rect 7904 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8072 7104
rect 8136 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8304 7104
rect 7904 6016 8304 7040
rect 7904 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8072 6016
rect 8136 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8304 6016
rect 7904 4928 8304 5952
rect 7904 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8072 4928
rect 8136 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8304 4928
rect 7904 3840 8304 4864
rect 7904 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8072 3840
rect 8136 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8304 3840
rect 7904 3294 8304 3776
rect 7904 3058 7986 3294
rect 8222 3058 8304 3294
rect 7904 2752 8304 3058
rect 7904 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8072 2752
rect 8136 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8304 2752
rect 7904 934 8304 2688
rect 7904 698 7986 934
rect 8222 698 8304 934
rect 7904 -4 8304 698
rect 8644 26618 9044 26660
rect 8644 26382 8726 26618
rect 8962 26382 9044 26618
rect 8644 23968 9044 26382
rect 8644 23904 8652 23968
rect 8716 23904 8732 23968
rect 8796 23904 8812 23968
rect 8876 23904 8892 23968
rect 8956 23904 8972 23968
rect 9036 23904 9044 23968
rect 8644 22880 9044 23904
rect 8644 22816 8652 22880
rect 8716 22816 8732 22880
rect 8796 22816 8812 22880
rect 8876 22816 8892 22880
rect 8956 22816 8972 22880
rect 9036 22816 9044 22880
rect 8644 22034 9044 22816
rect 8644 21798 8726 22034
rect 8962 21798 9044 22034
rect 8644 21792 9044 21798
rect 8644 21728 8652 21792
rect 8716 21728 8732 21792
rect 8796 21728 8812 21792
rect 8876 21728 8892 21792
rect 8956 21728 8972 21792
rect 9036 21728 9044 21792
rect 8644 20704 9044 21728
rect 8644 20640 8652 20704
rect 8716 20640 8732 20704
rect 8796 20640 8812 20704
rect 8876 20640 8892 20704
rect 8956 20640 8972 20704
rect 9036 20640 9044 20704
rect 8644 19616 9044 20640
rect 8644 19552 8652 19616
rect 8716 19552 8732 19616
rect 8796 19552 8812 19616
rect 8876 19552 8892 19616
rect 8956 19552 8972 19616
rect 9036 19552 9044 19616
rect 8644 18528 9044 19552
rect 8644 18464 8652 18528
rect 8716 18464 8732 18528
rect 8796 18464 8812 18528
rect 8876 18464 8892 18528
rect 8956 18464 8972 18528
rect 9036 18464 9044 18528
rect 8644 17440 9044 18464
rect 8644 17376 8652 17440
rect 8716 17376 8732 17440
rect 8796 17376 8812 17440
rect 8876 17376 8892 17440
rect 8956 17376 8972 17440
rect 9036 17376 9044 17440
rect 8644 16352 9044 17376
rect 8644 16288 8652 16352
rect 8716 16288 8732 16352
rect 8796 16288 8812 16352
rect 8876 16288 8892 16352
rect 8956 16288 8972 16352
rect 9036 16288 9044 16352
rect 8644 16034 9044 16288
rect 8644 15798 8726 16034
rect 8962 15798 9044 16034
rect 8644 15264 9044 15798
rect 8644 15200 8652 15264
rect 8716 15200 8732 15264
rect 8796 15200 8812 15264
rect 8876 15200 8892 15264
rect 8956 15200 8972 15264
rect 9036 15200 9044 15264
rect 8644 14176 9044 15200
rect 8644 14112 8652 14176
rect 8716 14112 8732 14176
rect 8796 14112 8812 14176
rect 8876 14112 8892 14176
rect 8956 14112 8972 14176
rect 9036 14112 9044 14176
rect 8644 13088 9044 14112
rect 8644 13024 8652 13088
rect 8716 13024 8732 13088
rect 8796 13024 8812 13088
rect 8876 13024 8892 13088
rect 8956 13024 8972 13088
rect 9036 13024 9044 13088
rect 8644 12000 9044 13024
rect 13904 25958 14304 26660
rect 13904 25722 13986 25958
rect 14222 25722 14304 25958
rect 13904 24512 14304 25722
rect 13904 24448 13912 24512
rect 13976 24448 13992 24512
rect 14056 24448 14072 24512
rect 14136 24448 14152 24512
rect 14216 24448 14232 24512
rect 14296 24448 14304 24512
rect 13904 23424 14304 24448
rect 13904 23360 13912 23424
rect 13976 23360 13992 23424
rect 14056 23360 14072 23424
rect 14136 23360 14152 23424
rect 14216 23360 14232 23424
rect 14296 23360 14304 23424
rect 13904 22336 14304 23360
rect 13904 22272 13912 22336
rect 13976 22272 13992 22336
rect 14056 22272 14072 22336
rect 14136 22272 14152 22336
rect 14216 22272 14232 22336
rect 14296 22272 14304 22336
rect 13904 21294 14304 22272
rect 13904 21248 13986 21294
rect 14222 21248 14304 21294
rect 13904 21184 13912 21248
rect 13976 21184 13986 21248
rect 14222 21184 14232 21248
rect 14296 21184 14304 21248
rect 13904 21058 13986 21184
rect 14222 21058 14304 21184
rect 13904 20160 14304 21058
rect 13904 20096 13912 20160
rect 13976 20096 13992 20160
rect 14056 20096 14072 20160
rect 14136 20096 14152 20160
rect 14216 20096 14232 20160
rect 14296 20096 14304 20160
rect 13904 19072 14304 20096
rect 13904 19008 13912 19072
rect 13976 19008 13992 19072
rect 14056 19008 14072 19072
rect 14136 19008 14152 19072
rect 14216 19008 14232 19072
rect 14296 19008 14304 19072
rect 13904 17984 14304 19008
rect 13904 17920 13912 17984
rect 13976 17920 13992 17984
rect 14056 17920 14072 17984
rect 14136 17920 14152 17984
rect 14216 17920 14232 17984
rect 14296 17920 14304 17984
rect 13904 16896 14304 17920
rect 13904 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14152 16896
rect 14216 16832 14232 16896
rect 14296 16832 14304 16896
rect 13904 15808 14304 16832
rect 13904 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14152 15808
rect 14216 15744 14232 15808
rect 14296 15744 14304 15808
rect 13904 15294 14304 15744
rect 13904 15058 13986 15294
rect 14222 15058 14304 15294
rect 13904 14720 14304 15058
rect 13904 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14152 14720
rect 14216 14656 14232 14720
rect 14296 14656 14304 14720
rect 13904 13632 14304 14656
rect 13904 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14152 13632
rect 14216 13568 14232 13632
rect 14296 13568 14304 13632
rect 9443 12748 9509 12749
rect 9443 12684 9444 12748
rect 9508 12684 9509 12748
rect 9443 12683 9509 12684
rect 8644 11936 8652 12000
rect 8716 11936 8732 12000
rect 8796 11936 8812 12000
rect 8876 11936 8892 12000
rect 8956 11936 8972 12000
rect 9036 11936 9044 12000
rect 8644 10912 9044 11936
rect 8644 10848 8652 10912
rect 8716 10848 8732 10912
rect 8796 10848 8812 10912
rect 8876 10848 8892 10912
rect 8956 10848 8972 10912
rect 9036 10848 9044 10912
rect 8644 10034 9044 10848
rect 9446 10709 9506 12683
rect 13904 12544 14304 13568
rect 13904 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14152 12544
rect 14216 12480 14232 12544
rect 14296 12480 14304 12544
rect 13904 11456 14304 12480
rect 13904 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14152 11456
rect 14216 11392 14232 11456
rect 14296 11392 14304 11456
rect 9443 10708 9509 10709
rect 9443 10644 9444 10708
rect 9508 10644 9509 10708
rect 9443 10643 9509 10644
rect 8644 9824 8726 10034
rect 8962 9824 9044 10034
rect 8644 9760 8652 9824
rect 8716 9798 8726 9824
rect 8962 9798 8972 9824
rect 8716 9760 8732 9798
rect 8796 9760 8812 9798
rect 8876 9760 8892 9798
rect 8956 9760 8972 9798
rect 9036 9760 9044 9824
rect 8644 8736 9044 9760
rect 8644 8672 8652 8736
rect 8716 8672 8732 8736
rect 8796 8672 8812 8736
rect 8876 8672 8892 8736
rect 8956 8672 8972 8736
rect 9036 8672 9044 8736
rect 8644 7648 9044 8672
rect 8644 7584 8652 7648
rect 8716 7584 8732 7648
rect 8796 7584 8812 7648
rect 8876 7584 8892 7648
rect 8956 7584 8972 7648
rect 9036 7584 9044 7648
rect 8644 6560 9044 7584
rect 8644 6496 8652 6560
rect 8716 6496 8732 6560
rect 8796 6496 8812 6560
rect 8876 6496 8892 6560
rect 8956 6496 8972 6560
rect 9036 6496 9044 6560
rect 8644 5472 9044 6496
rect 8644 5408 8652 5472
rect 8716 5408 8732 5472
rect 8796 5408 8812 5472
rect 8876 5408 8892 5472
rect 8956 5408 8972 5472
rect 9036 5408 9044 5472
rect 8644 4384 9044 5408
rect 8644 4320 8652 4384
rect 8716 4320 8732 4384
rect 8796 4320 8812 4384
rect 8876 4320 8892 4384
rect 8956 4320 8972 4384
rect 9036 4320 9044 4384
rect 8644 4034 9044 4320
rect 8644 3798 8726 4034
rect 8962 3798 9044 4034
rect 8644 3296 9044 3798
rect 8644 3232 8652 3296
rect 8716 3232 8732 3296
rect 8796 3232 8812 3296
rect 8876 3232 8892 3296
rect 8956 3232 8972 3296
rect 9036 3232 9044 3296
rect 8644 2208 9044 3232
rect 8644 2144 8652 2208
rect 8716 2144 8732 2208
rect 8796 2144 8812 2208
rect 8876 2144 8892 2208
rect 8956 2144 8972 2208
rect 9036 2144 9044 2208
rect 8644 274 9044 2144
rect 8644 38 8726 274
rect 8962 38 9044 274
rect 8644 -4 9044 38
rect 13904 10368 14304 11392
rect 13904 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14152 10368
rect 14216 10304 14232 10368
rect 14296 10304 14304 10368
rect 13904 9294 14304 10304
rect 13904 9280 13986 9294
rect 14222 9280 14304 9294
rect 13904 9216 13912 9280
rect 13976 9216 13986 9280
rect 14222 9216 14232 9280
rect 14296 9216 14304 9280
rect 13904 9058 13986 9216
rect 14222 9058 14304 9216
rect 13904 8192 14304 9058
rect 13904 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14152 8192
rect 14216 8128 14232 8192
rect 14296 8128 14304 8192
rect 13904 7104 14304 8128
rect 13904 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14152 7104
rect 14216 7040 14232 7104
rect 14296 7040 14304 7104
rect 13904 6016 14304 7040
rect 13904 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14152 6016
rect 14216 5952 14232 6016
rect 14296 5952 14304 6016
rect 13904 4928 14304 5952
rect 13904 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14152 4928
rect 14216 4864 14232 4928
rect 14296 4864 14304 4928
rect 13904 3840 14304 4864
rect 13904 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14152 3840
rect 14216 3776 14232 3840
rect 14296 3776 14304 3840
rect 13904 3294 14304 3776
rect 13904 3058 13986 3294
rect 14222 3058 14304 3294
rect 13904 2752 14304 3058
rect 13904 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14152 2752
rect 14216 2688 14232 2752
rect 14296 2688 14304 2752
rect 13904 934 14304 2688
rect 13904 698 13986 934
rect 14222 698 14304 934
rect 13904 -4 14304 698
rect 14644 26618 15044 26660
rect 14644 26382 14726 26618
rect 14962 26382 15044 26618
rect 14644 23968 15044 26382
rect 14644 23904 14652 23968
rect 14716 23904 14732 23968
rect 14796 23904 14812 23968
rect 14876 23904 14892 23968
rect 14956 23904 14972 23968
rect 15036 23904 15044 23968
rect 14644 22880 15044 23904
rect 14644 22816 14652 22880
rect 14716 22816 14732 22880
rect 14796 22816 14812 22880
rect 14876 22816 14892 22880
rect 14956 22816 14972 22880
rect 15036 22816 15044 22880
rect 14644 22034 15044 22816
rect 14644 21798 14726 22034
rect 14962 21798 15044 22034
rect 14644 21792 15044 21798
rect 14644 21728 14652 21792
rect 14716 21728 14732 21792
rect 14796 21728 14812 21792
rect 14876 21728 14892 21792
rect 14956 21728 14972 21792
rect 15036 21728 15044 21792
rect 14644 20704 15044 21728
rect 14644 20640 14652 20704
rect 14716 20640 14732 20704
rect 14796 20640 14812 20704
rect 14876 20640 14892 20704
rect 14956 20640 14972 20704
rect 15036 20640 15044 20704
rect 14644 19616 15044 20640
rect 14644 19552 14652 19616
rect 14716 19552 14732 19616
rect 14796 19552 14812 19616
rect 14876 19552 14892 19616
rect 14956 19552 14972 19616
rect 15036 19552 15044 19616
rect 14644 18528 15044 19552
rect 14644 18464 14652 18528
rect 14716 18464 14732 18528
rect 14796 18464 14812 18528
rect 14876 18464 14892 18528
rect 14956 18464 14972 18528
rect 15036 18464 15044 18528
rect 14644 17440 15044 18464
rect 14644 17376 14652 17440
rect 14716 17376 14732 17440
rect 14796 17376 14812 17440
rect 14876 17376 14892 17440
rect 14956 17376 14972 17440
rect 15036 17376 15044 17440
rect 14644 16352 15044 17376
rect 14644 16288 14652 16352
rect 14716 16288 14732 16352
rect 14796 16288 14812 16352
rect 14876 16288 14892 16352
rect 14956 16288 14972 16352
rect 15036 16288 15044 16352
rect 14644 16034 15044 16288
rect 14644 15798 14726 16034
rect 14962 15798 15044 16034
rect 14644 15264 15044 15798
rect 14644 15200 14652 15264
rect 14716 15200 14732 15264
rect 14796 15200 14812 15264
rect 14876 15200 14892 15264
rect 14956 15200 14972 15264
rect 15036 15200 15044 15264
rect 14644 14176 15044 15200
rect 14644 14112 14652 14176
rect 14716 14112 14732 14176
rect 14796 14112 14812 14176
rect 14876 14112 14892 14176
rect 14956 14112 14972 14176
rect 15036 14112 15044 14176
rect 14644 13088 15044 14112
rect 14644 13024 14652 13088
rect 14716 13024 14732 13088
rect 14796 13024 14812 13088
rect 14876 13024 14892 13088
rect 14956 13024 14972 13088
rect 15036 13024 15044 13088
rect 14644 12000 15044 13024
rect 14644 11936 14652 12000
rect 14716 11936 14732 12000
rect 14796 11936 14812 12000
rect 14876 11936 14892 12000
rect 14956 11936 14972 12000
rect 15036 11936 15044 12000
rect 14644 10912 15044 11936
rect 14644 10848 14652 10912
rect 14716 10848 14732 10912
rect 14796 10848 14812 10912
rect 14876 10848 14892 10912
rect 14956 10848 14972 10912
rect 15036 10848 15044 10912
rect 14644 10034 15044 10848
rect 14644 9824 14726 10034
rect 14962 9824 15044 10034
rect 14644 9760 14652 9824
rect 14716 9798 14726 9824
rect 14962 9798 14972 9824
rect 14716 9760 14732 9798
rect 14796 9760 14812 9798
rect 14876 9760 14892 9798
rect 14956 9760 14972 9798
rect 15036 9760 15044 9824
rect 14644 8736 15044 9760
rect 14644 8672 14652 8736
rect 14716 8672 14732 8736
rect 14796 8672 14812 8736
rect 14876 8672 14892 8736
rect 14956 8672 14972 8736
rect 15036 8672 15044 8736
rect 14644 7648 15044 8672
rect 14644 7584 14652 7648
rect 14716 7584 14732 7648
rect 14796 7584 14812 7648
rect 14876 7584 14892 7648
rect 14956 7584 14972 7648
rect 15036 7584 15044 7648
rect 14644 6560 15044 7584
rect 14644 6496 14652 6560
rect 14716 6496 14732 6560
rect 14796 6496 14812 6560
rect 14876 6496 14892 6560
rect 14956 6496 14972 6560
rect 15036 6496 15044 6560
rect 14644 5472 15044 6496
rect 14644 5408 14652 5472
rect 14716 5408 14732 5472
rect 14796 5408 14812 5472
rect 14876 5408 14892 5472
rect 14956 5408 14972 5472
rect 15036 5408 15044 5472
rect 14644 4384 15044 5408
rect 14644 4320 14652 4384
rect 14716 4320 14732 4384
rect 14796 4320 14812 4384
rect 14876 4320 14892 4384
rect 14956 4320 14972 4384
rect 15036 4320 15044 4384
rect 14644 4034 15044 4320
rect 14644 3798 14726 4034
rect 14962 3798 15044 4034
rect 14644 3296 15044 3798
rect 14644 3232 14652 3296
rect 14716 3232 14732 3296
rect 14796 3232 14812 3296
rect 14876 3232 14892 3296
rect 14956 3232 14972 3296
rect 15036 3232 15044 3296
rect 14644 2208 15044 3232
rect 14644 2144 14652 2208
rect 14716 2144 14732 2208
rect 14796 2144 14812 2208
rect 14876 2144 14892 2208
rect 14956 2144 14972 2208
rect 15036 2144 15044 2208
rect 14644 274 15044 2144
rect 14644 38 14726 274
rect 14962 38 15044 274
rect 14644 -4 15044 38
rect 19904 25958 20304 26660
rect 19904 25722 19986 25958
rect 20222 25722 20304 25958
rect 19904 24512 20304 25722
rect 19904 24448 19912 24512
rect 19976 24448 19992 24512
rect 20056 24448 20072 24512
rect 20136 24448 20152 24512
rect 20216 24448 20232 24512
rect 20296 24448 20304 24512
rect 19904 23424 20304 24448
rect 19904 23360 19912 23424
rect 19976 23360 19992 23424
rect 20056 23360 20072 23424
rect 20136 23360 20152 23424
rect 20216 23360 20232 23424
rect 20296 23360 20304 23424
rect 19904 22336 20304 23360
rect 19904 22272 19912 22336
rect 19976 22272 19992 22336
rect 20056 22272 20072 22336
rect 20136 22272 20152 22336
rect 20216 22272 20232 22336
rect 20296 22272 20304 22336
rect 19904 21294 20304 22272
rect 19904 21248 19986 21294
rect 20222 21248 20304 21294
rect 19904 21184 19912 21248
rect 19976 21184 19986 21248
rect 20222 21184 20232 21248
rect 20296 21184 20304 21248
rect 19904 21058 19986 21184
rect 20222 21058 20304 21184
rect 19904 20160 20304 21058
rect 19904 20096 19912 20160
rect 19976 20096 19992 20160
rect 20056 20096 20072 20160
rect 20136 20096 20152 20160
rect 20216 20096 20232 20160
rect 20296 20096 20304 20160
rect 19904 19072 20304 20096
rect 19904 19008 19912 19072
rect 19976 19008 19992 19072
rect 20056 19008 20072 19072
rect 20136 19008 20152 19072
rect 20216 19008 20232 19072
rect 20296 19008 20304 19072
rect 19904 17984 20304 19008
rect 19904 17920 19912 17984
rect 19976 17920 19992 17984
rect 20056 17920 20072 17984
rect 20136 17920 20152 17984
rect 20216 17920 20232 17984
rect 20296 17920 20304 17984
rect 19904 16896 20304 17920
rect 19904 16832 19912 16896
rect 19976 16832 19992 16896
rect 20056 16832 20072 16896
rect 20136 16832 20152 16896
rect 20216 16832 20232 16896
rect 20296 16832 20304 16896
rect 19904 15808 20304 16832
rect 19904 15744 19912 15808
rect 19976 15744 19992 15808
rect 20056 15744 20072 15808
rect 20136 15744 20152 15808
rect 20216 15744 20232 15808
rect 20296 15744 20304 15808
rect 19904 15294 20304 15744
rect 19904 15058 19986 15294
rect 20222 15058 20304 15294
rect 19904 14720 20304 15058
rect 19904 14656 19912 14720
rect 19976 14656 19992 14720
rect 20056 14656 20072 14720
rect 20136 14656 20152 14720
rect 20216 14656 20232 14720
rect 20296 14656 20304 14720
rect 19904 13632 20304 14656
rect 19904 13568 19912 13632
rect 19976 13568 19992 13632
rect 20056 13568 20072 13632
rect 20136 13568 20152 13632
rect 20216 13568 20232 13632
rect 20296 13568 20304 13632
rect 19904 12544 20304 13568
rect 19904 12480 19912 12544
rect 19976 12480 19992 12544
rect 20056 12480 20072 12544
rect 20136 12480 20152 12544
rect 20216 12480 20232 12544
rect 20296 12480 20304 12544
rect 19904 11456 20304 12480
rect 19904 11392 19912 11456
rect 19976 11392 19992 11456
rect 20056 11392 20072 11456
rect 20136 11392 20152 11456
rect 20216 11392 20232 11456
rect 20296 11392 20304 11456
rect 19904 10368 20304 11392
rect 19904 10304 19912 10368
rect 19976 10304 19992 10368
rect 20056 10304 20072 10368
rect 20136 10304 20152 10368
rect 20216 10304 20232 10368
rect 20296 10304 20304 10368
rect 19904 9294 20304 10304
rect 19904 9280 19986 9294
rect 20222 9280 20304 9294
rect 19904 9216 19912 9280
rect 19976 9216 19986 9280
rect 20222 9216 20232 9280
rect 20296 9216 20304 9280
rect 19904 9058 19986 9216
rect 20222 9058 20304 9216
rect 19904 8192 20304 9058
rect 19904 8128 19912 8192
rect 19976 8128 19992 8192
rect 20056 8128 20072 8192
rect 20136 8128 20152 8192
rect 20216 8128 20232 8192
rect 20296 8128 20304 8192
rect 19904 7104 20304 8128
rect 19904 7040 19912 7104
rect 19976 7040 19992 7104
rect 20056 7040 20072 7104
rect 20136 7040 20152 7104
rect 20216 7040 20232 7104
rect 20296 7040 20304 7104
rect 19904 6016 20304 7040
rect 19904 5952 19912 6016
rect 19976 5952 19992 6016
rect 20056 5952 20072 6016
rect 20136 5952 20152 6016
rect 20216 5952 20232 6016
rect 20296 5952 20304 6016
rect 19904 4928 20304 5952
rect 19904 4864 19912 4928
rect 19976 4864 19992 4928
rect 20056 4864 20072 4928
rect 20136 4864 20152 4928
rect 20216 4864 20232 4928
rect 20296 4864 20304 4928
rect 19904 3840 20304 4864
rect 19904 3776 19912 3840
rect 19976 3776 19992 3840
rect 20056 3776 20072 3840
rect 20136 3776 20152 3840
rect 20216 3776 20232 3840
rect 20296 3776 20304 3840
rect 19904 3294 20304 3776
rect 19904 3058 19986 3294
rect 20222 3058 20304 3294
rect 19904 2752 20304 3058
rect 19904 2688 19912 2752
rect 19976 2688 19992 2752
rect 20056 2688 20072 2752
rect 20136 2688 20152 2752
rect 20216 2688 20232 2752
rect 20296 2688 20304 2752
rect 19904 934 20304 2688
rect 19904 698 19986 934
rect 20222 698 20304 934
rect 19904 -4 20304 698
rect 20644 26618 21044 26660
rect 20644 26382 20726 26618
rect 20962 26382 21044 26618
rect 20644 23968 21044 26382
rect 25688 26618 26008 26660
rect 25688 26382 25730 26618
rect 25966 26382 26008 26618
rect 20644 23904 20652 23968
rect 20716 23904 20732 23968
rect 20796 23904 20812 23968
rect 20876 23904 20892 23968
rect 20956 23904 20972 23968
rect 21036 23904 21044 23968
rect 20644 22880 21044 23904
rect 20644 22816 20652 22880
rect 20716 22816 20732 22880
rect 20796 22816 20812 22880
rect 20876 22816 20892 22880
rect 20956 22816 20972 22880
rect 21036 22816 21044 22880
rect 20644 22034 21044 22816
rect 20644 21798 20726 22034
rect 20962 21798 21044 22034
rect 20644 21792 21044 21798
rect 20644 21728 20652 21792
rect 20716 21728 20732 21792
rect 20796 21728 20812 21792
rect 20876 21728 20892 21792
rect 20956 21728 20972 21792
rect 21036 21728 21044 21792
rect 20644 20704 21044 21728
rect 20644 20640 20652 20704
rect 20716 20640 20732 20704
rect 20796 20640 20812 20704
rect 20876 20640 20892 20704
rect 20956 20640 20972 20704
rect 21036 20640 21044 20704
rect 20644 19616 21044 20640
rect 20644 19552 20652 19616
rect 20716 19552 20732 19616
rect 20796 19552 20812 19616
rect 20876 19552 20892 19616
rect 20956 19552 20972 19616
rect 21036 19552 21044 19616
rect 20644 18528 21044 19552
rect 20644 18464 20652 18528
rect 20716 18464 20732 18528
rect 20796 18464 20812 18528
rect 20876 18464 20892 18528
rect 20956 18464 20972 18528
rect 21036 18464 21044 18528
rect 20644 17440 21044 18464
rect 20644 17376 20652 17440
rect 20716 17376 20732 17440
rect 20796 17376 20812 17440
rect 20876 17376 20892 17440
rect 20956 17376 20972 17440
rect 21036 17376 21044 17440
rect 20644 16352 21044 17376
rect 20644 16288 20652 16352
rect 20716 16288 20732 16352
rect 20796 16288 20812 16352
rect 20876 16288 20892 16352
rect 20956 16288 20972 16352
rect 21036 16288 21044 16352
rect 20644 16034 21044 16288
rect 20644 15798 20726 16034
rect 20962 15798 21044 16034
rect 20644 15264 21044 15798
rect 20644 15200 20652 15264
rect 20716 15200 20732 15264
rect 20796 15200 20812 15264
rect 20876 15200 20892 15264
rect 20956 15200 20972 15264
rect 21036 15200 21044 15264
rect 20644 14176 21044 15200
rect 20644 14112 20652 14176
rect 20716 14112 20732 14176
rect 20796 14112 20812 14176
rect 20876 14112 20892 14176
rect 20956 14112 20972 14176
rect 21036 14112 21044 14176
rect 20644 13088 21044 14112
rect 20644 13024 20652 13088
rect 20716 13024 20732 13088
rect 20796 13024 20812 13088
rect 20876 13024 20892 13088
rect 20956 13024 20972 13088
rect 21036 13024 21044 13088
rect 20644 12000 21044 13024
rect 20644 11936 20652 12000
rect 20716 11936 20732 12000
rect 20796 11936 20812 12000
rect 20876 11936 20892 12000
rect 20956 11936 20972 12000
rect 21036 11936 21044 12000
rect 20644 10912 21044 11936
rect 20644 10848 20652 10912
rect 20716 10848 20732 10912
rect 20796 10848 20812 10912
rect 20876 10848 20892 10912
rect 20956 10848 20972 10912
rect 21036 10848 21044 10912
rect 20644 10034 21044 10848
rect 20644 9824 20726 10034
rect 20962 9824 21044 10034
rect 20644 9760 20652 9824
rect 20716 9798 20726 9824
rect 20962 9798 20972 9824
rect 20716 9760 20732 9798
rect 20796 9760 20812 9798
rect 20876 9760 20892 9798
rect 20956 9760 20972 9798
rect 21036 9760 21044 9824
rect 20644 8736 21044 9760
rect 20644 8672 20652 8736
rect 20716 8672 20732 8736
rect 20796 8672 20812 8736
rect 20876 8672 20892 8736
rect 20956 8672 20972 8736
rect 21036 8672 21044 8736
rect 20644 7648 21044 8672
rect 20644 7584 20652 7648
rect 20716 7584 20732 7648
rect 20796 7584 20812 7648
rect 20876 7584 20892 7648
rect 20956 7584 20972 7648
rect 21036 7584 21044 7648
rect 20644 6560 21044 7584
rect 20644 6496 20652 6560
rect 20716 6496 20732 6560
rect 20796 6496 20812 6560
rect 20876 6496 20892 6560
rect 20956 6496 20972 6560
rect 21036 6496 21044 6560
rect 20644 5472 21044 6496
rect 20644 5408 20652 5472
rect 20716 5408 20732 5472
rect 20796 5408 20812 5472
rect 20876 5408 20892 5472
rect 20956 5408 20972 5472
rect 21036 5408 21044 5472
rect 20644 4384 21044 5408
rect 20644 4320 20652 4384
rect 20716 4320 20732 4384
rect 20796 4320 20812 4384
rect 20876 4320 20892 4384
rect 20956 4320 20972 4384
rect 21036 4320 21044 4384
rect 20644 4034 21044 4320
rect 20644 3798 20726 4034
rect 20962 3798 21044 4034
rect 20644 3296 21044 3798
rect 20644 3232 20652 3296
rect 20716 3232 20732 3296
rect 20796 3232 20812 3296
rect 20876 3232 20892 3296
rect 20956 3232 20972 3296
rect 21036 3232 21044 3296
rect 20644 2208 21044 3232
rect 20644 2144 20652 2208
rect 20716 2144 20732 2208
rect 20796 2144 20812 2208
rect 20876 2144 20892 2208
rect 20956 2144 20972 2208
rect 21036 2144 21044 2208
rect 20644 274 21044 2144
rect 25028 25958 25348 26000
rect 25028 25722 25070 25958
rect 25306 25722 25348 25958
rect 25028 21294 25348 25722
rect 25028 21058 25070 21294
rect 25306 21058 25348 21294
rect 25028 15294 25348 21058
rect 25028 15058 25070 15294
rect 25306 15058 25348 15294
rect 25028 9294 25348 15058
rect 25028 9058 25070 9294
rect 25306 9058 25348 9294
rect 25028 3294 25348 9058
rect 25028 3058 25070 3294
rect 25306 3058 25348 3294
rect 25028 934 25348 3058
rect 25028 698 25070 934
rect 25306 698 25348 934
rect 25028 656 25348 698
rect 25688 22034 26008 26382
rect 25688 21798 25730 22034
rect 25966 21798 26008 22034
rect 25688 16034 26008 21798
rect 25688 15798 25730 16034
rect 25966 15798 26008 16034
rect 25688 10034 26008 15798
rect 25688 9798 25730 10034
rect 25966 9798 26008 10034
rect 25688 4034 26008 9798
rect 25688 3798 25730 4034
rect 25966 3798 26008 4034
rect 20644 38 20726 274
rect 20962 38 21044 274
rect 20644 -4 21044 38
rect 25688 274 26008 3798
rect 25688 38 25730 274
rect 25966 38 26008 274
rect 25688 -4 26008 38
<< via4 >>
rect -1034 26382 -798 26618
rect -1034 21798 -798 22034
rect -1034 15798 -798 16034
rect -1034 9798 -798 10034
rect -1034 3798 -798 4034
rect -374 25722 -138 25958
rect -374 21058 -138 21294
rect -374 15058 -138 15294
rect -374 9058 -138 9294
rect -374 3058 -138 3294
rect -374 698 -138 934
rect 1986 25722 2222 25958
rect 1986 21248 2222 21294
rect 1986 21184 1992 21248
rect 1992 21184 2056 21248
rect 2056 21184 2072 21248
rect 2072 21184 2136 21248
rect 2136 21184 2152 21248
rect 2152 21184 2216 21248
rect 2216 21184 2222 21248
rect 1986 21058 2222 21184
rect 1986 15058 2222 15294
rect 1986 9280 2222 9294
rect 1986 9216 1992 9280
rect 1992 9216 2056 9280
rect 2056 9216 2072 9280
rect 2072 9216 2136 9280
rect 2136 9216 2152 9280
rect 2152 9216 2216 9280
rect 2216 9216 2222 9280
rect 1986 9058 2222 9216
rect 1986 3058 2222 3294
rect 1986 698 2222 934
rect -1034 38 -798 274
rect 2726 26382 2962 26618
rect 2726 21798 2962 22034
rect 2726 15798 2962 16034
rect 2726 9824 2962 10034
rect 2726 9798 2732 9824
rect 2732 9798 2796 9824
rect 2796 9798 2812 9824
rect 2812 9798 2876 9824
rect 2876 9798 2892 9824
rect 2892 9798 2956 9824
rect 2956 9798 2962 9824
rect 2726 3798 2962 4034
rect 2726 38 2962 274
rect 7986 25722 8222 25958
rect 7986 21248 8222 21294
rect 7986 21184 7992 21248
rect 7992 21184 8056 21248
rect 8056 21184 8072 21248
rect 8072 21184 8136 21248
rect 8136 21184 8152 21248
rect 8152 21184 8216 21248
rect 8216 21184 8222 21248
rect 7986 21058 8222 21184
rect 7986 15058 8222 15294
rect 7986 9280 8222 9294
rect 7986 9216 7992 9280
rect 7992 9216 8056 9280
rect 8056 9216 8072 9280
rect 8072 9216 8136 9280
rect 8136 9216 8152 9280
rect 8152 9216 8216 9280
rect 8216 9216 8222 9280
rect 7986 9058 8222 9216
rect 7986 3058 8222 3294
rect 7986 698 8222 934
rect 8726 26382 8962 26618
rect 8726 21798 8962 22034
rect 8726 15798 8962 16034
rect 13986 25722 14222 25958
rect 13986 21248 14222 21294
rect 13986 21184 13992 21248
rect 13992 21184 14056 21248
rect 14056 21184 14072 21248
rect 14072 21184 14136 21248
rect 14136 21184 14152 21248
rect 14152 21184 14216 21248
rect 14216 21184 14222 21248
rect 13986 21058 14222 21184
rect 13986 15058 14222 15294
rect 8726 9824 8962 10034
rect 8726 9798 8732 9824
rect 8732 9798 8796 9824
rect 8796 9798 8812 9824
rect 8812 9798 8876 9824
rect 8876 9798 8892 9824
rect 8892 9798 8956 9824
rect 8956 9798 8962 9824
rect 8726 3798 8962 4034
rect 8726 38 8962 274
rect 13986 9280 14222 9294
rect 13986 9216 13992 9280
rect 13992 9216 14056 9280
rect 14056 9216 14072 9280
rect 14072 9216 14136 9280
rect 14136 9216 14152 9280
rect 14152 9216 14216 9280
rect 14216 9216 14222 9280
rect 13986 9058 14222 9216
rect 13986 3058 14222 3294
rect 13986 698 14222 934
rect 14726 26382 14962 26618
rect 14726 21798 14962 22034
rect 14726 15798 14962 16034
rect 14726 9824 14962 10034
rect 14726 9798 14732 9824
rect 14732 9798 14796 9824
rect 14796 9798 14812 9824
rect 14812 9798 14876 9824
rect 14876 9798 14892 9824
rect 14892 9798 14956 9824
rect 14956 9798 14962 9824
rect 14726 3798 14962 4034
rect 14726 38 14962 274
rect 19986 25722 20222 25958
rect 19986 21248 20222 21294
rect 19986 21184 19992 21248
rect 19992 21184 20056 21248
rect 20056 21184 20072 21248
rect 20072 21184 20136 21248
rect 20136 21184 20152 21248
rect 20152 21184 20216 21248
rect 20216 21184 20222 21248
rect 19986 21058 20222 21184
rect 19986 15058 20222 15294
rect 19986 9280 20222 9294
rect 19986 9216 19992 9280
rect 19992 9216 20056 9280
rect 20056 9216 20072 9280
rect 20072 9216 20136 9280
rect 20136 9216 20152 9280
rect 20152 9216 20216 9280
rect 20216 9216 20222 9280
rect 19986 9058 20222 9216
rect 19986 3058 20222 3294
rect 19986 698 20222 934
rect 20726 26382 20962 26618
rect 25730 26382 25966 26618
rect 20726 21798 20962 22034
rect 20726 15798 20962 16034
rect 20726 9824 20962 10034
rect 20726 9798 20732 9824
rect 20732 9798 20796 9824
rect 20796 9798 20812 9824
rect 20812 9798 20876 9824
rect 20876 9798 20892 9824
rect 20892 9798 20956 9824
rect 20956 9798 20962 9824
rect 20726 3798 20962 4034
rect 25070 25722 25306 25958
rect 25070 21058 25306 21294
rect 25070 15058 25306 15294
rect 25070 9058 25306 9294
rect 25070 3058 25306 3294
rect 25070 698 25306 934
rect 25730 21798 25966 22034
rect 25730 15798 25966 16034
rect 25730 9798 25966 10034
rect 25730 3798 25966 4034
rect 20726 38 20962 274
rect 25730 38 25966 274
<< metal5 >>
rect -1076 26618 26008 26660
rect -1076 26382 -1034 26618
rect -798 26382 2726 26618
rect 2962 26382 8726 26618
rect 8962 26382 14726 26618
rect 14962 26382 20726 26618
rect 20962 26382 25730 26618
rect 25966 26382 26008 26618
rect -1076 26340 26008 26382
rect -416 25958 25348 26000
rect -416 25722 -374 25958
rect -138 25722 1986 25958
rect 2222 25722 7986 25958
rect 8222 25722 13986 25958
rect 14222 25722 19986 25958
rect 20222 25722 25070 25958
rect 25306 25722 25348 25958
rect -416 25680 25348 25722
rect -1076 22034 26008 22116
rect -1076 21798 -1034 22034
rect -798 21798 2726 22034
rect 2962 21798 8726 22034
rect 8962 21798 14726 22034
rect 14962 21798 20726 22034
rect 20962 21798 25730 22034
rect 25966 21798 26008 22034
rect -1076 21716 26008 21798
rect -1076 21294 26008 21376
rect -1076 21058 -374 21294
rect -138 21058 1986 21294
rect 2222 21058 7986 21294
rect 8222 21058 13986 21294
rect 14222 21058 19986 21294
rect 20222 21058 25070 21294
rect 25306 21058 26008 21294
rect -1076 20976 26008 21058
rect -1076 16034 26008 16116
rect -1076 15798 -1034 16034
rect -798 15798 2726 16034
rect 2962 15798 8726 16034
rect 8962 15798 14726 16034
rect 14962 15798 20726 16034
rect 20962 15798 25730 16034
rect 25966 15798 26008 16034
rect -1076 15716 26008 15798
rect -1076 15294 26008 15376
rect -1076 15058 -374 15294
rect -138 15058 1986 15294
rect 2222 15058 7986 15294
rect 8222 15058 13986 15294
rect 14222 15058 19986 15294
rect 20222 15058 25070 15294
rect 25306 15058 26008 15294
rect -1076 14976 26008 15058
rect -1076 10034 26008 10116
rect -1076 9798 -1034 10034
rect -798 9798 2726 10034
rect 2962 9798 8726 10034
rect 8962 9798 14726 10034
rect 14962 9798 20726 10034
rect 20962 9798 25730 10034
rect 25966 9798 26008 10034
rect -1076 9716 26008 9798
rect -1076 9294 26008 9376
rect -1076 9058 -374 9294
rect -138 9058 1986 9294
rect 2222 9058 7986 9294
rect 8222 9058 13986 9294
rect 14222 9058 19986 9294
rect 20222 9058 25070 9294
rect 25306 9058 26008 9294
rect -1076 8976 26008 9058
rect -1076 4034 26008 4116
rect -1076 3798 -1034 4034
rect -798 3798 2726 4034
rect 2962 3798 8726 4034
rect 8962 3798 14726 4034
rect 14962 3798 20726 4034
rect 20962 3798 25730 4034
rect 25966 3798 26008 4034
rect -1076 3716 26008 3798
rect -1076 3294 26008 3376
rect -1076 3058 -374 3294
rect -138 3058 1986 3294
rect 2222 3058 7986 3294
rect 8222 3058 13986 3294
rect 14222 3058 19986 3294
rect 20222 3058 25070 3294
rect 25306 3058 26008 3294
rect -1076 2976 26008 3058
rect -416 934 25348 976
rect -416 698 -374 934
rect -138 698 1986 934
rect 2222 698 7986 934
rect 8222 698 13986 934
rect 14222 698 19986 934
rect 20222 698 25070 934
rect 25306 698 25348 934
rect -416 656 25348 698
rect -1076 274 26008 316
rect -1076 38 -1034 274
rect -798 38 2726 274
rect 2962 38 8726 274
rect 8962 38 14726 274
rect 14962 38 20726 274
rect 20962 38 25730 274
rect 25966 38 26008 274
rect -1076 -4 26008 38
use sky130_fd_sc_hd__buf_2  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12052 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _246_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 17204 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 14260 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _248_
timestamp 1701704242
transform -1 0 14628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _249_
timestamp 1701704242
transform 1 0 15088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _250_
timestamp 1701704242
transform 1 0 17388 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _251_
timestamp 1701704242
transform -1 0 18400 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _252_
timestamp 1701704242
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _253_
timestamp 1701704242
transform 1 0 18492 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _254_
timestamp 1701704242
transform -1 0 19136 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _255_
timestamp 1701704242
transform 1 0 21068 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _256_
timestamp 1701704242
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _257_
timestamp 1701704242
transform 1 0 23276 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _258_
timestamp 1701704242
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _259_
timestamp 1701704242
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _260_
timestamp 1701704242
transform 1 0 13892 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _261_
timestamp 1701704242
transform 1 0 21344 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _262_
timestamp 1701704242
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _263_
timestamp 1701704242
transform 1 0 18584 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _264_
timestamp 1701704242
transform -1 0 19044 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _265_
timestamp 1701704242
transform -1 0 16928 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _266_
timestamp 1701704242
transform -1 0 11408 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _267_
timestamp 1701704242
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _268_
timestamp 1701704242
transform -1 0 14628 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _269_
timestamp 1701704242
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _270_
timestamp 1701704242
transform -1 0 14536 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _271_
timestamp 1701704242
transform -1 0 12052 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _272_
timestamp 1701704242
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _273_
timestamp 1701704242
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _274_
timestamp 1701704242
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _275_
timestamp 1701704242
transform 1 0 16008 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _276_
timestamp 1701704242
transform 1 0 11040 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _277_
timestamp 1701704242
transform -1 0 14536 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _278_
timestamp 1701704242
transform 1 0 12144 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _279_
timestamp 1701704242
transform -1 0 10212 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _280_
timestamp 1701704242
transform -1 0 4784 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _281_
timestamp 1701704242
transform -1 0 12052 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _282_
timestamp 1701704242
transform 1 0 4508 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _283_
timestamp 1701704242
transform -1 0 10672 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _284_
timestamp 1701704242
transform -1 0 1748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _285_
timestamp 1701704242
transform -1 0 12052 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _286_
timestamp 1701704242
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _287_
timestamp 1701704242
transform -1 0 11868 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _288_
timestamp 1701704242
transform -1 0 8832 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _289_
timestamp 1701704242
transform 1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _290_
timestamp 1701704242
transform -1 0 9476 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _291_
timestamp 1701704242
transform 1 0 3220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _292_
timestamp 1701704242
transform -1 0 12052 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _293_
timestamp 1701704242
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _294_
timestamp 1701704242
transform -1 0 8740 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _295_
timestamp 1701704242
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _296_
timestamp 1701704242
transform -1 0 6992 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _297_
timestamp 1701704242
transform -1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _298_
timestamp 1701704242
transform -1 0 9476 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _299_
timestamp 1701704242
transform -1 0 2392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _300_
timestamp 1701704242
transform -1 0 9476 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _301_
timestamp 1701704242
transform 1 0 3128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _302_
timestamp 1701704242
transform -1 0 9568 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _303_
timestamp 1701704242
transform -1 0 1840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _304_
timestamp 1701704242
transform -1 0 9568 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _305_
timestamp 1701704242
transform -1 0 7360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _306_
timestamp 1701704242
transform 1 0 9016 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _307_
timestamp 1701704242
transform 1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _308_
timestamp 1701704242
transform 1 0 10856 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _309_
timestamp 1701704242
transform 1 0 10396 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _310_
timestamp 1701704242
transform 1 0 11592 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _311_
timestamp 1701704242
transform 1 0 11500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _312_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 15640 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _313_
timestamp 1701704242
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _314_
timestamp 1701704242
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315__61 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 14352 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316__62
timestamp 1701704242
transform 1 0 5888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317__63
timestamp 1701704242
transform 1 0 6348 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318__64
timestamp 1701704242
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319__65
timestamp 1701704242
transform 1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320__66
timestamp 1701704242
transform 1 0 2484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321__67
timestamp 1701704242
transform 1 0 1840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322__68
timestamp 1701704242
transform -1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323__69
timestamp 1701704242
transform -1 0 2208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324__70
timestamp 1701704242
transform -1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _325_
timestamp 1701704242
transform -1 0 11776 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326__71
timestamp 1701704242
transform -1 0 2668 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327__72
timestamp 1701704242
transform -1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328__73
timestamp 1701704242
transform -1 0 6992 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329__74
timestamp 1701704242
transform -1 0 1840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330__75
timestamp 1701704242
transform -1 0 4232 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331__76
timestamp 1701704242
transform 1 0 4232 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332__77
timestamp 1701704242
transform 1 0 9292 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333__78
timestamp 1701704242
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334__79
timestamp 1701704242
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335__80
timestamp 1701704242
transform 1 0 9292 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _336_
timestamp 1701704242
transform 1 0 13616 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337__81
timestamp 1701704242
transform -1 0 18308 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338__82
timestamp 1701704242
transform -1 0 18584 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339__83
timestamp 1701704242
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340__84
timestamp 1701704242
transform -1 0 19044 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341__85
timestamp 1701704242
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342__86
timestamp 1701704242
transform -1 0 16928 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343__87
timestamp 1701704242
transform 1 0 21344 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344__88
timestamp 1701704242
transform -1 0 15824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345__89
timestamp 1701704242
transform -1 0 18952 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346__90
timestamp 1701704242
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _347_
timestamp 1701704242
transform -1 0 14904 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348__91
timestamp 1701704242
transform -1 0 14352 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349__92
timestamp 1701704242
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350__93
timestamp 1701704242
transform 1 0 10396 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351__94
timestamp 1701704242
transform -1 0 6900 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352__95
timestamp 1701704242
transform -1 0 12052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353__96
timestamp 1701704242
transform -1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354__97
timestamp 1701704242
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355__98
timestamp 1701704242
transform 1 0 2760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356__99
timestamp 1701704242
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357__100
timestamp 1701704242
transform -1 0 1840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _358_
timestamp 1701704242
transform 1 0 1564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359__101
timestamp 1701704242
transform -1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360__102
timestamp 1701704242
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361__103
timestamp 1701704242
transform 1 0 2668 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362__104
timestamp 1701704242
transform 1 0 2668 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363__105
timestamp 1701704242
transform 1 0 8464 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364__106
timestamp 1701704242
transform 1 0 12144 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365__107
timestamp 1701704242
transform -1 0 4508 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366__108
timestamp 1701704242
transform 1 0 6440 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367__109
timestamp 1701704242
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368__110
timestamp 1701704242
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _369_
timestamp 1701704242
transform 1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370__111
timestamp 1701704242
transform -1 0 13984 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371__112
timestamp 1701704242
transform -1 0 11040 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372__113
timestamp 1701704242
transform -1 0 18952 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373__114
timestamp 1701704242
transform -1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374__115
timestamp 1701704242
transform -1 0 21620 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375__116
timestamp 1701704242
transform 1 0 21068 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376__117
timestamp 1701704242
transform -1 0 21712 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377__118
timestamp 1701704242
transform -1 0 21528 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378__119
timestamp 1701704242
transform 1 0 23276 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379__120
timestamp 1701704242
transform -1 0 16376 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _380_
timestamp 1701704242
transform 1 0 2208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _381__121
timestamp 1701704242
transform 1 0 23276 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _382__122
timestamp 1701704242
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _383__123
timestamp 1701704242
transform -1 0 16468 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _384__124
timestamp 1701704242
transform -1 0 15824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _385__125
timestamp 1701704242
transform 1 0 16192 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386__126
timestamp 1701704242
transform -1 0 14536 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _387__127
timestamp 1701704242
transform -1 0 12604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388__128
timestamp 1701704242
transform -1 0 13524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _389__129
timestamp 1701704242
transform -1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _390__130
timestamp 1701704242
transform -1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _391_
timestamp 1701704242
transform -1 0 11500 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _392__131
timestamp 1701704242
transform -1 0 8464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _393__132
timestamp 1701704242
transform -1 0 9200 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _394__133
timestamp 1701704242
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _395__134
timestamp 1701704242
transform -1 0 1840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _396__135
timestamp 1701704242
transform -1 0 4140 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _397__136
timestamp 1701704242
transform -1 0 4048 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _398__137
timestamp 1701704242
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _399__138
timestamp 1701704242
transform 1 0 13432 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _400__139
timestamp 1701704242
transform -1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _401__140
timestamp 1701704242
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _402_
timestamp 1701704242
transform 1 0 13616 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _403__141
timestamp 1701704242
transform -1 0 14352 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _404__142
timestamp 1701704242
transform -1 0 9568 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _405__143
timestamp 1701704242
transform -1 0 13248 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _406__144
timestamp 1701704242
transform -1 0 13800 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _407__145
timestamp 1701704242
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _408__146
timestamp 1701704242
transform 1 0 17940 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _409__147
timestamp 1701704242
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _410__148
timestamp 1701704242
transform 1 0 16192 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _411__149
timestamp 1701704242
transform 1 0 23276 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _412__150
timestamp 1701704242
transform 1 0 23276 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _413_
timestamp 1701704242
transform 1 0 6440 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _414__151
timestamp 1701704242
transform -1 0 21620 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _415__152
timestamp 1701704242
transform 1 0 23276 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _416__153
timestamp 1701704242
transform -1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _417__154
timestamp 1701704242
transform -1 0 21712 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _418__155
timestamp 1701704242
transform -1 0 18952 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _419__156
timestamp 1701704242
transform -1 0 17020 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _420__157
timestamp 1701704242
transform -1 0 13248 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _421__158
timestamp 1701704242
transform -1 0 14076 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _422__159
timestamp 1701704242
transform -1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _423__160
timestamp 1701704242
transform -1 0 13248 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _424_
timestamp 1701704242
transform 1 0 2300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _425__1
timestamp 1701704242
transform 1 0 4048 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _426__2
timestamp 1701704242
transform 1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _427__3
timestamp 1701704242
transform -1 0 2668 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _428__4
timestamp 1701704242
transform -1 0 6716 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _429__5
timestamp 1701704242
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _430__6
timestamp 1701704242
transform 1 0 1564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _431__7
timestamp 1701704242
transform 1 0 3956 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _432__8
timestamp 1701704242
transform 1 0 1564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433__9
timestamp 1701704242
transform 1 0 6440 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _434__10
timestamp 1701704242
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _435_
timestamp 1701704242
transform 1 0 1564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _436__11
timestamp 1701704242
transform -1 0 9200 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _437__12
timestamp 1701704242
transform -1 0 8832 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _438__13
timestamp 1701704242
transform -1 0 14444 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _439__14
timestamp 1701704242
transform 1 0 14352 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _440__15
timestamp 1701704242
transform 1 0 9660 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _441__16
timestamp 1701704242
transform 1 0 11592 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _442__17
timestamp 1701704242
transform 1 0 20516 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _443__18
timestamp 1701704242
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _444__19
timestamp 1701704242
transform 1 0 19320 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _445__20
timestamp 1701704242
transform -1 0 14352 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _446_
timestamp 1701704242
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _447__21
timestamp 1701704242
transform 1 0 21252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _448__22
timestamp 1701704242
transform -1 0 22080 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _449__23
timestamp 1701704242
transform -1 0 23368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450__24
timestamp 1701704242
transform 1 0 23276 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _451__25
timestamp 1701704242
transform -1 0 21528 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _452__26
timestamp 1701704242
transform 1 0 23276 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _453__27
timestamp 1701704242
transform -1 0 16928 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _454__28
timestamp 1701704242
transform -1 0 19136 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _455__29
timestamp 1701704242
transform -1 0 14536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _456__30
timestamp 1701704242
transform -1 0 13616 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _457_
timestamp 1701704242
transform -1 0 9292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _458__31
timestamp 1701704242
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _459__32
timestamp 1701704242
transform -1 0 7728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _460__33
timestamp 1701704242
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _461__34
timestamp 1701704242
transform 1 0 6440 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _462__35
timestamp 1701704242
transform -1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _463__36
timestamp 1701704242
transform 1 0 12052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _464__37
timestamp 1701704242
transform 1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _465__38
timestamp 1701704242
transform -1 0 6992 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _466__39
timestamp 1701704242
transform 1 0 4140 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _467__40
timestamp 1701704242
transform -1 0 3772 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _468_
timestamp 1701704242
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _469__41
timestamp 1701704242
transform 1 0 9016 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _470__42
timestamp 1701704242
transform -1 0 6716 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _471__43
timestamp 1701704242
transform 1 0 6716 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _472__44
timestamp 1701704242
transform -1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _473__45
timestamp 1701704242
transform 1 0 15180 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _474__46
timestamp 1701704242
transform -1 0 15548 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _475__47
timestamp 1701704242
transform -1 0 13984 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _476__48
timestamp 1701704242
transform -1 0 14536 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _477__49
timestamp 1701704242
transform 1 0 18584 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _478__50
timestamp 1701704242
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _479_
timestamp 1701704242
transform 1 0 14352 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _480__51
timestamp 1701704242
transform -1 0 21620 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _481__52
timestamp 1701704242
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _482__53
timestamp 1701704242
transform -1 0 22908 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _483__54
timestamp 1701704242
transform 1 0 23276 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _484__55
timestamp 1701704242
transform -1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _485__56
timestamp 1701704242
transform 1 0 23092 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _486__57
timestamp 1701704242
transform 1 0 23276 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _487__58
timestamp 1701704242
transform 1 0 23276 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _488__59
timestamp 1701704242
transform -1 0 16560 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _489__60
timestamp 1701704242
transform -1 0 21344 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 11408 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _491_
timestamp 1701704242
transform 1 0 6348 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _492_
timestamp 1701704242
transform 1 0 8464 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _493_
timestamp 1701704242
transform 1 0 7360 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _494_
timestamp 1701704242
transform 1 0 2208 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _495_
timestamp 1701704242
transform -1 0 3312 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _496_
timestamp 1701704242
transform 1 0 3312 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _497_
timestamp 1701704242
transform 1 0 5520 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _498_
timestamp 1701704242
transform 1 0 1748 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _499_
timestamp 1701704242
transform 1 0 2208 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _500_
timestamp 1701704242
transform 1 0 1840 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _501_
timestamp 1701704242
transform 1 0 1840 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _502_
timestamp 1701704242
transform -1 0 6440 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _503_
timestamp 1701704242
transform 1 0 4784 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _504_
timestamp 1701704242
transform 1 0 3864 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _505_
timestamp 1701704242
transform 1 0 4508 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _506_
timestamp 1701704242
transform 1 0 9568 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _507_
timestamp 1701704242
transform -1 0 11040 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _508_
timestamp 1701704242
transform -1 0 11408 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _509_
timestamp 1701704242
transform 1 0 10580 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _510_
timestamp 1701704242
transform 1 0 14996 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _511_
timestamp 1701704242
transform 1 0 14720 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _512_
timestamp 1701704242
transform 1 0 17664 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _513_
timestamp 1701704242
transform -1 0 15916 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _514_
timestamp 1701704242
transform -1 0 20700 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _515_
timestamp 1701704242
transform 1 0 17296 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _516_
timestamp 1701704242
transform -1 0 20332 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _517_
timestamp 1701704242
transform -1 0 15548 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _518_
timestamp 1701704242
transform -1 0 18952 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _519_
timestamp 1701704242
transform -1 0 19964 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _520_
timestamp 1701704242
transform -1 0 13984 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _521_
timestamp 1701704242
transform -1 0 13984 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _522_
timestamp 1701704242
transform 1 0 10764 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _523_
timestamp 1701704242
transform 1 0 11592 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _524_
timestamp 1701704242
transform -1 0 11408 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _525_
timestamp 1701704242
transform 1 0 9292 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _526_
timestamp 1701704242
transform 1 0 4324 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _527_
timestamp 1701704242
transform 1 0 3312 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _528_
timestamp 1701704242
transform 1 0 2208 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _529_
timestamp 1701704242
transform 1 0 9200 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _530_
timestamp 1701704242
transform 1 0 1840 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _531_
timestamp 1701704242
transform 1 0 3312 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _532_
timestamp 1701704242
transform 1 0 4784 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _533_
timestamp 1701704242
transform 1 0 3864 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _534_
timestamp 1701704242
transform -1 0 8832 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _535_
timestamp 1701704242
transform -1 0 8832 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _536_
timestamp 1701704242
transform 1 0 5336 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _537_
timestamp 1701704242
transform -1 0 6808 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _538_
timestamp 1701704242
transform 1 0 11040 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _539_
timestamp 1701704242
transform 1 0 11040 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _540_
timestamp 1701704242
transform 1 0 12052 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _541_
timestamp 1701704242
transform 1 0 11868 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _542_
timestamp 1701704242
transform -1 0 18308 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _543_
timestamp 1701704242
transform -1 0 18584 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _544_
timestamp 1701704242
transform -1 0 19136 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _545_
timestamp 1701704242
transform -1 0 18492 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _546_
timestamp 1701704242
transform 1 0 20700 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _547_
timestamp 1701704242
transform 1 0 19228 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _548_
timestamp 1701704242
transform -1 0 23092 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _549_
timestamp 1701704242
transform 1 0 14904 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _550_
timestamp 1701704242
transform -1 0 21252 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _551_
timestamp 1701704242
transform 1 0 19596 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _552_
timestamp 1701704242
transform 1 0 16008 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _553_
timestamp 1701704242
transform 1 0 14996 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _554_
timestamp 1701704242
transform 1 0 10672 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _555_
timestamp 1701704242
transform -1 0 13616 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _556_
timestamp 1701704242
transform 1 0 9936 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _557_
timestamp 1701704242
transform -1 0 12972 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _558_
timestamp 1701704242
transform 1 0 4324 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _559_
timestamp 1701704242
transform 1 0 3312 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _560_
timestamp 1701704242
transform -1 0 6256 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _561_
timestamp 1701704242
transform -1 0 10396 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _562_
timestamp 1701704242
transform 1 0 4784 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _563_
timestamp 1701704242
transform 1 0 3312 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _564_
timestamp 1701704242
transform -1 0 6256 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _565_
timestamp 1701704242
transform 1 0 4784 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _566_
timestamp 1701704242
transform -1 0 9568 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _567_
timestamp 1701704242
transform 1 0 7636 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _568_
timestamp 1701704242
transform 1 0 6808 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _569_
timestamp 1701704242
transform 1 0 6532 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _570_
timestamp 1701704242
transform 1 0 12512 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _571_
timestamp 1701704242
transform 1 0 11500 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _572_
timestamp 1701704242
transform -1 0 13524 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _573_
timestamp 1701704242
transform -1 0 13524 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _574_
timestamp 1701704242
transform 1 0 18308 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _575_
timestamp 1701704242
transform 1 0 17388 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _576_
timestamp 1701704242
transform -1 0 21160 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _577_
timestamp 1701704242
transform -1 0 15824 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _578_
timestamp 1701704242
transform 1 0 21804 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _579_
timestamp 1701704242
transform 1 0 21804 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _580_
timestamp 1701704242
transform -1 0 21436 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _581_
timestamp 1701704242
transform -1 0 17112 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _582_
timestamp 1701704242
transform 1 0 21804 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _583_
timestamp 1701704242
transform 1 0 21804 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _584_
timestamp 1701704242
transform -1 0 17020 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _585_
timestamp 1701704242
transform -1 0 19596 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _586_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 15640 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _587_
timestamp 1701704242
transform -1 0 14260 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _588_
timestamp 1701704242
transform 1 0 11040 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _589_
timestamp 1701704242
transform -1 0 12972 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _590_
timestamp 1701704242
transform 1 0 4048 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _591_
timestamp 1701704242
transform 1 0 4324 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _592_
timestamp 1701704242
transform 1 0 3220 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _593_
timestamp 1701704242
transform -1 0 7360 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _594_
timestamp 1701704242
transform 1 0 4324 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _595_
timestamp 1701704242
transform 1 0 4416 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _596_
timestamp 1701704242
transform -1 0 4784 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _597_
timestamp 1701704242
transform 1 0 4416 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _598_
timestamp 1701704242
transform 1 0 9568 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _599_
timestamp 1701704242
transform -1 0 7912 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _600_
timestamp 1701704242
transform 1 0 6808 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _601_
timestamp 1701704242
transform 1 0 6624 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _602_
timestamp 1701704242
transform -1 0 13984 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _603_
timestamp 1701704242
transform 1 0 12512 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _604_
timestamp 1701704242
transform 1 0 14076 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _605_
timestamp 1701704242
transform 1 0 13340 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _606_
timestamp 1701704242
transform 1 0 19228 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _607_
timestamp 1701704242
transform 1 0 18860 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _608_
timestamp 1701704242
transform 1 0 19964 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _609_
timestamp 1701704242
transform 1 0 16652 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _610_
timestamp 1701704242
transform -1 0 21436 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _611_
timestamp 1701704242
transform -1 0 22172 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _612_
timestamp 1701704242
transform 1 0 20700 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _613_
timestamp 1701704242
transform 1 0 18492 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _614_
timestamp 1701704242
transform 1 0 19228 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _615_
timestamp 1701704242
transform -1 0 20424 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _616_
timestamp 1701704242
transform -1 0 18492 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _617_
timestamp 1701704242
transform 1 0 16652 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _618_
timestamp 1701704242
transform 1 0 12144 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _619_
timestamp 1701704242
transform 1 0 12512 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _620_
timestamp 1701704242
transform -1 0 13800 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _621_
timestamp 1701704242
transform -1 0 13800 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _622_
timestamp 1701704242
transform 1 0 6348 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _623_
timestamp 1701704242
transform 1 0 4784 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _624_
timestamp 1701704242
transform -1 0 5520 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _625_
timestamp 1701704242
transform -1 0 6256 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _626_
timestamp 1701704242
transform -1 0 6256 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _627_
timestamp 1701704242
transform 1 0 4048 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _628_
timestamp 1701704242
transform 1 0 4784 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _629_
timestamp 1701704242
transform -1 0 6808 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _630_
timestamp 1701704242
transform -1 0 8188 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _631_
timestamp 1701704242
transform 1 0 9660 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _632_
timestamp 1701704242
transform -1 0 8464 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _633_
timestamp 1701704242
transform -1 0 8464 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _634_
timestamp 1701704242
transform 1 0 14076 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _635_
timestamp 1701704242
transform 1 0 12972 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _636_
timestamp 1701704242
transform 1 0 12052 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _637_
timestamp 1701704242
transform 1 0 12052 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _638_
timestamp 1701704242
transform 1 0 19596 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _639_
timestamp 1701704242
transform 1 0 19228 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _640_
timestamp 1701704242
transform 1 0 19596 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _641_
timestamp 1701704242
transform 1 0 15548 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _642_
timestamp 1701704242
transform 1 0 21804 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _643_
timestamp 1701704242
transform -1 0 23276 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _644_
timestamp 1701704242
transform 1 0 20700 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _645_
timestamp 1701704242
transform -1 0 19780 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _646_
timestamp 1701704242
transform 1 0 20700 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _647_
timestamp 1701704242
transform -1 0 23276 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _648_
timestamp 1701704242
transform -1 0 16100 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _649_
timestamp 1701704242
transform -1 0 18124 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _650_
timestamp 1701704242
transform 1 0 9568 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _651_
timestamp 1701704242
transform 1 0 7360 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _652_
timestamp 1701704242
transform 1 0 6992 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _653_
timestamp 1701704242
transform -1 0 11040 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _654_
timestamp 1701704242
transform 1 0 1840 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _655_
timestamp 1701704242
transform 1 0 2208 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _656_
timestamp 1701704242
transform -1 0 4784 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _657_
timestamp 1701704242
transform 1 0 8464 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _658_
timestamp 1701704242
transform -1 0 3312 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _659_
timestamp 1701704242
transform -1 0 3680 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _660_
timestamp 1701704242
transform 1 0 3312 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _661_
timestamp 1701704242
transform 1 0 3312 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _662_
timestamp 1701704242
transform 1 0 6624 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _663_
timestamp 1701704242
transform -1 0 10488 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _664_
timestamp 1701704242
transform 1 0 4784 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _665_
timestamp 1701704242
transform 1 0 4784 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _666_
timestamp 1701704242
transform 1 0 10672 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _667_
timestamp 1701704242
transform 1 0 9936 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _668_
timestamp 1701704242
transform 1 0 9660 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _669_
timestamp 1701704242
transform 1 0 11776 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _670_
timestamp 1701704242
transform -1 0 19596 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _671_
timestamp 1701704242
transform 1 0 16652 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _672_
timestamp 1701704242
transform -1 0 19964 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _673_
timestamp 1701704242
transform 1 0 14720 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _674_
timestamp 1701704242
transform 1 0 16836 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _675_
timestamp 1701704242
transform -1 0 21252 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _676_
timestamp 1701704242
transform 1 0 19228 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _677_
timestamp 1701704242
transform 1 0 14076 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _678_
timestamp 1701704242
transform 1 0 19228 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _679_
timestamp 1701704242
transform 1 0 17204 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _680_
timestamp 1701704242
transform 1 0 14076 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _681_
timestamp 1701704242
transform 1 0 14076 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _682_
timestamp 1701704242
transform -1 0 13984 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _683_
timestamp 1701704242
transform -1 0 13800 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _684_
timestamp 1701704242
transform 1 0 8280 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _685_
timestamp 1701704242
transform -1 0 7268 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _686_
timestamp 1701704242
transform 1 0 7268 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _687_
timestamp 1701704242
transform 1 0 6992 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _688_
timestamp 1701704242
transform 1 0 4784 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _689_
timestamp 1701704242
transform 1 0 7360 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _690_
timestamp 1701704242
transform 1 0 4784 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _691_
timestamp 1701704242
transform 1 0 5520 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _692_
timestamp 1701704242
transform 1 0 5888 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _693_
timestamp 1701704242
transform 1 0 6348 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _694_
timestamp 1701704242
transform 1 0 9936 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _695_
timestamp 1701704242
transform 1 0 9936 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _696_
timestamp 1701704242
transform 1 0 8464 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _697_
timestamp 1701704242
transform 1 0 8096 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _698_
timestamp 1701704242
transform 1 0 15548 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _699_
timestamp 1701704242
transform 1 0 14444 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _700_
timestamp 1701704242
transform -1 0 13800 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _701_
timestamp 1701704242
transform -1 0 13800 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _702_
timestamp 1701704242
transform -1 0 17940 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _703_
timestamp 1701704242
transform 1 0 14536 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _704_
timestamp 1701704242
transform -1 0 20608 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _705_
timestamp 1701704242
transform 1 0 18124 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _706_
timestamp 1701704242
transform -1 0 23276 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _707_
timestamp 1701704242
transform -1 0 22540 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _708_
timestamp 1701704242
transform -1 0 21620 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _709_
timestamp 1701704242
transform -1 0 18584 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _710_
timestamp 1701704242
transform -1 0 23276 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _711_
timestamp 1701704242
transform -1 0 23092 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _712_
timestamp 1701704242
transform -1 0 16008 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _713_
timestamp 1701704242
transform -1 0 16192 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 12972 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__228_
timestamp 1701704242
transform 1 0 11500 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__229_
timestamp 1701704242
transform 1 0 6348 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__230_
timestamp 1701704242
transform -1 0 9292 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__231_
timestamp 1701704242
transform 1 0 15456 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__232_
timestamp 1701704242
transform -1 0 10580 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__233_
timestamp 1701704242
transform 1 0 8188 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__234_
timestamp 1701704242
transform 1 0 15824 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__235_
timestamp 1701704242
transform 1 0 12420 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__236_
timestamp 1701704242
transform -1 0 9660 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__237_
timestamp 1701704242
transform 1 0 16652 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__238_
timestamp 1701704242
transform 1 0 16652 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__239_
timestamp 1701704242
transform 1 0 7820 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__240_
timestamp 1701704242
transform 1 0 13984 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__241_
timestamp 1701704242
transform 1 0 17296 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__242_
timestamp 1701704242
transform 1 0 8924 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__243_
timestamp 1701704242
transform 1 0 12144 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__244_
timestamp 1701704242
transform 1 0 19228 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1701704242
transform 1 0 11592 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__227_
timestamp 1701704242
transform -1 0 10764 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__228_
timestamp 1701704242
transform -1 0 10948 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__229_
timestamp 1701704242
transform -1 0 5796 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__230_
timestamp 1701704242
transform -1 0 6624 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__231_
timestamp 1701704242
transform 1 0 16008 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__232_
timestamp 1701704242
transform -1 0 8188 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__233_
timestamp 1701704242
transform -1 0 8648 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__234_
timestamp 1701704242
transform -1 0 15732 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__235_
timestamp 1701704242
transform -1 0 11408 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__236_
timestamp 1701704242
transform 1 0 8924 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__237_
timestamp 1701704242
transform 1 0 18768 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__238_
timestamp 1701704242
transform -1 0 15916 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__239_
timestamp 1701704242
transform -1 0 8556 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__240_
timestamp 1701704242
transform -1 0 13892 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__241_
timestamp 1701704242
transform -1 0 16652 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__242_
timestamp 1701704242
transform -1 0 8832 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__243_
timestamp 1701704242
transform -1 0 11408 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__244_
timestamp 1701704242
transform -1 0 18492 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__227_
timestamp 1701704242
transform 1 0 13524 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__228_
timestamp 1701704242
transform 1 0 13064 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__229_
timestamp 1701704242
transform 1 0 8556 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__230_
timestamp 1701704242
transform 1 0 9568 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__231_
timestamp 1701704242
transform 1 0 15916 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__232_
timestamp 1701704242
transform 1 0 10672 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__233_
timestamp 1701704242
transform 1 0 8924 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__234_
timestamp 1701704242
transform 1 0 19228 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__235_
timestamp 1701704242
transform 1 0 15916 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__236_
timestamp 1701704242
transform -1 0 8832 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__237_
timestamp 1701704242
transform -1 0 17112 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__238_
timestamp 1701704242
transform 1 0 17940 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__239_
timestamp 1701704242
transform 1 0 7912 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__240_
timestamp 1701704242
transform 1 0 16192 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__241_
timestamp 1701704242
transform 1 0 19780 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__242_
timestamp 1701704242
transform -1 0 8832 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__243_
timestamp 1701704242
transform 1 0 14628 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__244_
timestamp 1701704242
transform 1 0 21160 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1701704242
transform -1 0 8004 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1701704242
transform 1 0 9476 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1701704242
transform -1 0 8280 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1701704242
transform -1 0 11408 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1701704242
transform -1 0 16468 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1701704242
transform 1 0 17020 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1701704242
transform -1 0 15916 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1701704242
transform 1 0 16928 0 -1 16320
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1701704242
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1701704242
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1701704242
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_63
timestamp 1701704242
transform 1 0 6900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1701704242
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_97 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1701704242
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_113
timestamp 1701704242
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_126
timestamp 1701704242
transform 1 0 12696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_135
timestamp 1701704242
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1701704242
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_150
timestamp 1701704242
transform 1 0 14904 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_162
timestamp 1701704242
transform 1 0 16008 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_169
timestamp 1701704242
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_182
timestamp 1701704242
transform 1 0 17848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_194
timestamp 1701704242
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1701704242
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1701704242
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1701704242
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1701704242
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_237
timestamp 1701704242
transform 1 0 22908 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_243
timestamp 1701704242
transform 1 0 23460 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1701704242
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1701704242
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1701704242
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1701704242
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1701704242
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1701704242
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1701704242
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1701704242
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1701704242
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1701704242
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1701704242
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1701704242
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_122
timestamp 1701704242
transform 1 0 12328 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_134
timestamp 1701704242
transform 1 0 13432 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_146
timestamp 1701704242
transform 1 0 14536 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_158 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 15640 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_166
timestamp 1701704242
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1701704242
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1701704242
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1701704242
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1701704242
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1701704242
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1701704242
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1701704242
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_237
timestamp 1701704242
transform 1 0 22908 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_243
timestamp 1701704242
transform 1 0 23460 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1701704242
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1701704242
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1701704242
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1701704242
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1701704242
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1701704242
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_65
timestamp 1701704242
transform 1 0 7084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_72
timestamp 1701704242
transform 1 0 7728 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_80
timestamp 1701704242
transform 1 0 8464 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_85
timestamp 1701704242
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_103
timestamp 1701704242
transform 1 0 10580 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_111
timestamp 1701704242
transform 1 0 11316 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_125
timestamp 1701704242
transform 1 0 12604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_137
timestamp 1701704242
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1701704242
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1701704242
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1701704242
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1701704242
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1701704242
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1701704242
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1701704242
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1701704242
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1701704242
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_233
timestamp 1701704242
transform 1 0 22540 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_241
timestamp 1701704242
transform 1 0 23276 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1701704242
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1701704242
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1701704242
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1701704242
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1701704242
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1701704242
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_57
timestamp 1701704242
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_61
timestamp 1701704242
transform 1 0 6716 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_76
timestamp 1701704242
transform 1 0 8096 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_80
timestamp 1701704242
transform 1 0 8464 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_132
timestamp 1701704242
transform 1 0 13248 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_144
timestamp 1701704242
transform 1 0 14352 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_156
timestamp 1701704242
transform 1 0 15456 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1701704242
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1701704242
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1701704242
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1701704242
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1701704242
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1701704242
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_225
timestamp 1701704242
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_241
timestamp 1701704242
transform 1 0 23276 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1701704242
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1701704242
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1701704242
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1701704242
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_41
timestamp 1701704242
transform 1 0 4876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_49
timestamp 1701704242
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_56
timestamp 1701704242
transform 1 0 6256 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 1701704242
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_108
timestamp 1701704242
transform 1 0 11040 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_135
timestamp 1701704242
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1701704242
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_141
timestamp 1701704242
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_146
timestamp 1701704242
transform 1 0 14536 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_158
timestamp 1701704242
transform 1 0 15640 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_173
timestamp 1701704242
transform 1 0 17020 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_185
timestamp 1701704242
transform 1 0 18124 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1701704242
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1701704242
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1701704242
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_221
timestamp 1701704242
transform 1 0 21436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_232
timestamp 1701704242
transform 1 0 22448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_3
timestamp 1701704242
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_12
timestamp 1701704242
transform 1 0 2208 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_20
timestamp 1701704242
transform 1 0 2944 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_25
timestamp 1701704242
transform 1 0 3404 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_31
timestamp 1701704242
transform 1 0 3956 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_51
timestamp 1701704242
transform 1 0 5796 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_73
timestamp 1701704242
transform 1 0 7820 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_77
timestamp 1701704242
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_94
timestamp 1701704242
transform 1 0 9752 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_113
timestamp 1701704242
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_121
timestamp 1701704242
transform 1 0 12236 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_155
timestamp 1701704242
transform 1 0 15364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_160
timestamp 1701704242
transform 1 0 15824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1701704242
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_188
timestamp 1701704242
transform 1 0 18400 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_194
timestamp 1701704242
transform 1 0 18952 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_206
timestamp 1701704242
transform 1 0 20056 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_218
timestamp 1701704242
transform 1 0 21160 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_222
timestamp 1701704242
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_225
timestamp 1701704242
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_237
timestamp 1701704242
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_3
timestamp 1701704242
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_14
timestamp 1701704242
transform 1 0 2392 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_24
timestamp 1701704242
transform 1 0 3312 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_67
timestamp 1701704242
transform 1 0 7268 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_85
timestamp 1701704242
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_121
timestamp 1701704242
transform 1 0 12236 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 1701704242
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_150
timestamp 1701704242
transform 1 0 14904 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_167
timestamp 1701704242
transform 1 0 16468 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_3
timestamp 1701704242
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_57
timestamp 1701704242
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_121
timestamp 1701704242
transform 1 0 12236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_140
timestamp 1701704242
transform 1 0 13984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_172
timestamp 1701704242
transform 1 0 16928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_192
timestamp 1701704242
transform 1 0 18768 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_12
timestamp 1701704242
transform 1 0 2208 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_52
timestamp 1701704242
transform 1 0 5888 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_64
timestamp 1701704242
transform 1 0 6992 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1701704242
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp 1701704242
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_125
timestamp 1701704242
transform 1 0 12604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_137
timestamp 1701704242
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_173
timestamp 1701704242
transform 1 0 17020 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_194
timestamp 1701704242
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_229
timestamp 1701704242
transform 1 0 22172 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_3
timestamp 1701704242
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_8
timestamp 1701704242
transform 1 0 1840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_12
timestamp 1701704242
transform 1 0 2208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_57
timestamp 1701704242
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_113
timestamp 1701704242
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_147
timestamp 1701704242
transform 1 0 14628 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1701704242
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1701704242
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_3
timestamp 1701704242
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_64
timestamp 1701704242
transform 1 0 6992 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_123
timestamp 1701704242
transform 1 0 12420 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_144
timestamp 1701704242
transform 1 0 14352 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 1701704242
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_205
timestamp 1701704242
transform 1 0 19964 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_242
timestamp 1701704242
transform 1 0 23368 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_3
timestamp 1701704242
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_91
timestamp 1701704242
transform 1 0 9476 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_113
timestamp 1701704242
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_146
timestamp 1701704242
transform 1 0 14536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1701704242
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_222
timestamp 1701704242
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_3
timestamp 1701704242
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_49
timestamp 1701704242
transform 1 0 5612 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_61
timestamp 1701704242
transform 1 0 6716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1701704242
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_229
timestamp 1701704242
transform 1 0 22172 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_3
timestamp 1701704242
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_15
timestamp 1701704242
transform 1 0 2484 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1701704242
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_117
timestamp 1701704242
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_146
timestamp 1701704242
transform 1 0 14536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1701704242
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_3
timestamp 1701704242
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_29
timestamp 1701704242
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_51
timestamp 1701704242
transform 1 0 5796 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_75
timestamp 1701704242
transform 1 0 8004 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_123
timestamp 1701704242
transform 1 0 12420 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_3
timestamp 1701704242
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_57
timestamp 1701704242
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_113
timestamp 1701704242
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_172
timestamp 1701704242
transform 1 0 16928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1701704242
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_3
timestamp 1701704242
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_29
timestamp 1701704242
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_35
timestamp 1701704242
transform 1 0 4324 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_62
timestamp 1701704242
transform 1 0 6808 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_105
timestamp 1701704242
transform 1 0 10764 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1701704242
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_175
timestamp 1701704242
transform 1 0 17204 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_242
timestamp 1701704242
transform 1 0 23368 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_3
timestamp 1701704242
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_113
timestamp 1701704242
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1701704242
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_29
timestamp 1701704242
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1701704242
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_160
timestamp 1701704242
transform 1 0 15824 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_217
timestamp 1701704242
transform 1 0 21068 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_238
timestamp 1701704242
transform 1 0 23000 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_3
timestamp 1701704242
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_107
timestamp 1701704242
transform 1 0 10948 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1701704242
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_169
timestamp 1701704242
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_222
timestamp 1701704242
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_113
timestamp 1701704242
transform 1 0 11500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_147
timestamp 1701704242
transform 1 0 14628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1701704242
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1701704242
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_94
timestamp 1701704242
transform 1 0 9752 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_158
timestamp 1701704242
transform 1 0 15640 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1701704242
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_29
timestamp 1701704242
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 1701704242
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1701704242
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_237
timestamp 1701704242
transform 1 0 22908 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_3
timestamp 1701704242
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_113
timestamp 1701704242
transform 1 0 11500 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_138
timestamp 1701704242
transform 1 0 13800 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1701704242
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1701704242
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_3
timestamp 1701704242
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_29
timestamp 1701704242
transform 1 0 3772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_85
timestamp 1701704242
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_102
timestamp 1701704242
transform 1 0 10488 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_135
timestamp 1701704242
transform 1 0 13524 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_9
timestamp 1701704242
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_57
timestamp 1701704242
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_97
timestamp 1701704242
transform 1 0 10028 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_146
timestamp 1701704242
transform 1 0 14536 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1701704242
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1701704242
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_3
timestamp 1701704242
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_12
timestamp 1701704242
transform 1 0 2208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_16
timestamp 1701704242
transform 1 0 2576 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_29
timestamp 1701704242
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_91
timestamp 1701704242
transform 1 0 9476 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_112
timestamp 1701704242
transform 1 0 11408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1701704242
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1701704242
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_200
timestamp 1701704242
transform 1 0 19504 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_237
timestamp 1701704242
transform 1 0 22908 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_9
timestamp 1701704242
transform 1 0 1932 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_21
timestamp 1701704242
transform 1 0 3036 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_57
timestamp 1701704242
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_116
timestamp 1701704242
transform 1 0 11776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_149
timestamp 1701704242
transform 1 0 14812 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1701704242
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_221
timestamp 1701704242
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1701704242
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_237
timestamp 1701704242
transform 1 0 22908 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1701704242
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1701704242
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1701704242
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_29
timestamp 1701704242
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_60
timestamp 1701704242
transform 1 0 6624 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_112
timestamp 1701704242
transform 1 0 11408 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_138
timestamp 1701704242
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_147
timestamp 1701704242
transform 1 0 14628 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_197
timestamp 1701704242
transform 1 0 19228 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_201
timestamp 1701704242
transform 1 0 19596 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_213
timestamp 1701704242
transform 1 0 20700 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_225
timestamp 1701704242
transform 1 0 21804 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_237
timestamp 1701704242
transform 1 0 22908 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_243
timestamp 1701704242
transform 1 0 23460 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1701704242
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1701704242
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_27
timestamp 1701704242
transform 1 0 3588 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_119
timestamp 1701704242
transform 1 0 12052 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1701704242
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1701704242
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1701704242
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_237
timestamp 1701704242
transform 1 0 22908 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_243
timestamp 1701704242
transform 1 0 23460 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1701704242
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1701704242
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1701704242
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_29
timestamp 1701704242
transform 1 0 3772 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_79
timestamp 1701704242
transform 1 0 8372 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1701704242
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1701704242
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_233
timestamp 1701704242
transform 1 0 22540 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_237
timestamp 1701704242
transform 1 0 22908 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1701704242
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1701704242
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_27
timestamp 1701704242
transform 1 0 3588 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_35
timestamp 1701704242
transform 1 0 4324 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_108
timestamp 1701704242
transform 1 0 11040 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_113
timestamp 1701704242
transform 1 0 11500 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_117
timestamp 1701704242
transform 1 0 11868 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_139
timestamp 1701704242
transform 1 0 13892 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_169
timestamp 1701704242
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_214
timestamp 1701704242
transform 1 0 20792 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_222
timestamp 1701704242
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1701704242
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_237
timestamp 1701704242
transform 1 0 22908 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1701704242
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1701704242
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1701704242
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_29
timestamp 1701704242
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_37
timestamp 1701704242
transform 1 0 4508 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_62
timestamp 1701704242
transform 1 0 6808 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1701704242
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_85
timestamp 1701704242
transform 1 0 8924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_141
timestamp 1701704242
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_213
timestamp 1701704242
transform 1 0 20700 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_225
timestamp 1701704242
transform 1 0 21804 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_237
timestamp 1701704242
transform 1 0 22908 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_243
timestamp 1701704242
transform 1 0 23460 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1701704242
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1701704242
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1701704242
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_39
timestamp 1701704242
transform 1 0 4692 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_57
timestamp 1701704242
transform 1 0 6348 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_161
timestamp 1701704242
transform 1 0 15916 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_209
timestamp 1701704242
transform 1 0 20332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1701704242
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1701704242
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_237
timestamp 1701704242
transform 1 0 22908 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_243
timestamp 1701704242
transform 1 0 23460 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1701704242
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1701704242
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1701704242
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_29
timestamp 1701704242
transform 1 0 3772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_33
timestamp 1701704242
transform 1 0 4140 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_53
timestamp 1701704242
transform 1 0 5980 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_88
timestamp 1701704242
transform 1 0 9200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_181
timestamp 1701704242
transform 1 0 17756 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_194
timestamp 1701704242
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_200
timestamp 1701704242
transform 1 0 19504 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_212
timestamp 1701704242
transform 1 0 20608 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_224
timestamp 1701704242
transform 1 0 21712 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_236
timestamp 1701704242
transform 1 0 22816 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1701704242
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1701704242
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1701704242
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1701704242
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1701704242
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1701704242
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_57
timestamp 1701704242
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_91
timestamp 1701704242
transform 1 0 9476 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_140
timestamp 1701704242
transform 1 0 13984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_145
timestamp 1701704242
transform 1 0 14444 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_157
timestamp 1701704242
transform 1 0 15548 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_166
timestamp 1701704242
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_177
timestamp 1701704242
transform 1 0 17388 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 1701704242
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 1701704242
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 1701704242
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1701704242
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1701704242
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_237
timestamp 1701704242
transform 1 0 22908 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_243
timestamp 1701704242
transform 1 0 23460 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1701704242
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1701704242
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1701704242
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1701704242
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1701704242
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1701704242
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1701704242
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_77
timestamp 1701704242
transform 1 0 8188 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_85
timestamp 1701704242
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_99
timestamp 1701704242
transform 1 0 10212 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_103
timestamp 1701704242
transform 1 0 10580 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_123
timestamp 1701704242
transform 1 0 12420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1701704242
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1701704242
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_147
timestamp 1701704242
transform 1 0 14628 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_156
timestamp 1701704242
transform 1 0 15456 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_168
timestamp 1701704242
transform 1 0 16560 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_180
timestamp 1701704242
transform 1 0 17664 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_192
timestamp 1701704242
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1701704242
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 1701704242
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 1701704242
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_233
timestamp 1701704242
transform 1 0 22540 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_241
timestamp 1701704242
transform 1 0 23276 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1701704242
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1701704242
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1701704242
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1701704242
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1701704242
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1701704242
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1701704242
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1701704242
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1701704242
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 1701704242
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_105
timestamp 1701704242
transform 1 0 10764 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1701704242
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1701704242
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1701704242
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 1701704242
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 1701704242
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 1701704242
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1701704242
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1701704242
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 1701704242
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 1701704242
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 1701704242
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 1701704242
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1701704242
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1701704242
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_237
timestamp 1701704242
transform 1 0 22908 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_243
timestamp 1701704242
transform 1 0 23460 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1701704242
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1701704242
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1701704242
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1701704242
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1701704242
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1701704242
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1701704242
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1701704242
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1701704242
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1701704242
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1701704242
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 1701704242
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 1701704242
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 1701704242
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1701704242
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1701704242
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 1701704242
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 1701704242
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_177
timestamp 1701704242
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 1701704242
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1701704242
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1701704242
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 1701704242
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 1701704242
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_233
timestamp 1701704242
transform 1 0 22540 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_241
timestamp 1701704242
transform 1 0 23276 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1701704242
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1701704242
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1701704242
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1701704242
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1701704242
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1701704242
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1701704242
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1701704242
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1701704242
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 1701704242
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 1701704242
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1701704242
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1701704242
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1701704242
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 1701704242
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 1701704242
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1701704242
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1701704242
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1701704242
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1701704242
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 1701704242
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 1701704242
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 1701704242
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1701704242
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1701704242
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_237
timestamp 1701704242
transform 1 0 22908 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_243
timestamp 1701704242
transform 1 0 23460 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1701704242
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1701704242
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1701704242
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1701704242
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1701704242
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_53
timestamp 1701704242
transform 1 0 5980 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_57
timestamp 1701704242
transform 1 0 6348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_69
timestamp 1701704242
transform 1 0 7452 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_79
timestamp 1701704242
transform 1 0 8372 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1701704242
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_94
timestamp 1701704242
transform 1 0 9752 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_106
timestamp 1701704242
transform 1 0 10856 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_122
timestamp 1701704242
transform 1 0 12328 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_134
timestamp 1701704242
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_162
timestamp 1701704242
transform 1 0 16008 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_169
timestamp 1701704242
transform 1 0 16652 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_181
timestamp 1701704242
transform 1 0 17756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_193
timestamp 1701704242
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1701704242
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1701704242
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_221
timestamp 1701704242
transform 1 0 21436 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_225
timestamp 1701704242
transform 1 0 21804 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_237
timestamp 1701704242
transform 1 0 22908 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_243
timestamp 1701704242
transform 1 0 23460 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 12328 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1701704242
transform -1 0 16468 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1701704242
transform -1 0 10304 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1701704242
transform -1 0 10396 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1701704242
transform -1 0 12696 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1701704242
transform -1 0 12052 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1701704242
transform -1 0 16284 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1701704242
transform 1 0 11684 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1701704242
transform 1 0 11040 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1701704242
transform -1 0 7452 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1701704242
transform -1 0 12328 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1701704242
transform 1 0 9200 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1701704242
transform 1 0 7360 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1701704242
transform -1 0 8832 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1701704242
transform -1 0 17388 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1701704242
transform -1 0 15272 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1701704242
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1701704242
transform 1 0 17848 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1701704242
transform -1 0 11408 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1701704242
transform -1 0 9660 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1701704242
transform -1 0 12328 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1701704242
transform -1 0 12144 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1701704242
transform -1 0 18676 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1701704242
transform 1 0 4232 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1701704242
transform -1 0 11132 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1701704242
transform -1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1701704242
transform -1 0 17388 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1701704242
transform -1 0 18492 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1701704242
transform -1 0 12236 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1701704242
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1701704242
transform -1 0 17756 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1701704242
transform 1 0 10396 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1701704242
transform 1 0 8924 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1701704242
transform -1 0 22724 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1701704242
transform 1 0 8188 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1701704242
transform -1 0 21160 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1701704242
transform 1 0 15548 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1701704242
transform -1 0 21344 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1701704242
transform -1 0 21344 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1701704242
transform -1 0 11316 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1701704242
transform 1 0 9660 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1701704242
transform -1 0 20976 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1701704242
transform 1 0 6900 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1701704242
transform -1 0 21068 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1701704242
transform 1 0 1472 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1701704242
transform -1 0 8832 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1701704242
transform 1 0 11776 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1701704242
transform -1 0 23552 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1701704242
transform 1 0 22540 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1701704242
transform 1 0 12604 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1701704242
transform -1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1701704242
transform -1 0 22448 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1701704242
transform -1 0 19964 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1701704242
transform -1 0 22908 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1701704242
transform 1 0 22080 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1701704242
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1701704242
transform -1 0 17388 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1701704242
transform -1 0 11500 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1701704242
transform -1 0 16560 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1701704242
transform 1 0 14720 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1701704242
transform -1 0 18860 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1701704242
transform -1 0 17664 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1701704242
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1701704242
transform -1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1701704242
transform 1 0 2576 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1701704242
transform 1 0 1472 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1701704242
transform 1 0 1472 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1701704242
transform 1 0 13248 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1701704242
transform 1 0 6624 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1701704242
transform 1 0 6072 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1701704242
transform 1 0 17756 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1701704242
transform -1 0 23276 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1701704242
transform 1 0 2576 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1701704242
transform -1 0 14812 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1701704242
transform 1 0 2208 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1701704242
transform -1 0 22632 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1701704242
transform -1 0 18124 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1701704242
transform -1 0 21436 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1701704242
transform 1 0 4600 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1701704242
transform -1 0 20240 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1701704242
transform -1 0 21712 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1701704242
transform -1 0 14536 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1701704242
transform 1 0 1472 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1701704242
transform 1 0 18124 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1701704242
transform -1 0 14260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1701704242
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1701704242
transform -1 0 11500 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1701704242
transform 1 0 18216 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1701704242
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1701704242
transform 1 0 13248 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1701704242
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1701704242
transform 1 0 14536 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1701704242
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1701704242
transform 1 0 4048 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1701704242
transform -1 0 22908 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1701704242
transform -1 0 20516 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1701704242
transform -1 0 21896 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1701704242
transform 1 0 2576 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1701704242
transform 1 0 4048 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1701704242
transform 1 0 2944 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1701704242
transform 1 0 1472 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1701704242
transform 1 0 13616 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1701704242
transform 1 0 8004 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1701704242
transform -1 0 9476 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10396 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_6  output2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 12696 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  output3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 1932 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output4
timestamp 1701704242
transform -1 0 1932 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  output5
timestamp 1701704242
transform 1 0 11500 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output6
timestamp 1701704242
transform -1 0 2208 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output7
timestamp 1701704242
transform 1 0 8924 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  output8
timestamp 1701704242
transform 1 0 7820 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output9
timestamp 1701704242
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output10
timestamp 1701704242
transform 1 0 14628 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  output11
timestamp 1701704242
transform 1 0 22724 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output12
timestamp 1701704242
transform 1 0 15180 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output13
timestamp 1701704242
transform 1 0 22724 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  output14
timestamp 1701704242
transform 1 0 23000 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output15
timestamp 1701704242
transform 1 0 23000 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output16
timestamp 1701704242
transform 1 0 23000 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output17
timestamp 1701704242
transform 1 0 23000 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output18
timestamp 1701704242
transform 1 0 22172 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output19
timestamp 1701704242
transform 1 0 23000 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output20
timestamp 1701704242
transform 1 0 22172 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  output21
timestamp 1701704242
transform 1 0 22724 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output22
timestamp 1701704242
transform 1 0 22724 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output23
timestamp 1701704242
transform 1 0 22724 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output24
timestamp 1701704242
transform 1 0 14076 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output25
timestamp 1701704242
transform -1 0 17848 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output26
timestamp 1701704242
transform 1 0 18124 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  output27
timestamp 1701704242
transform 1 0 12972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  output28
timestamp 1701704242
transform 1 0 6992 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output29
timestamp 1701704242
transform 1 0 7820 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output30
timestamp 1701704242
transform 1 0 5980 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output31
timestamp 1701704242
transform 1 0 11500 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output32
timestamp 1701704242
transform -1 0 2208 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output33
timestamp 1701704242
transform -1 0 2208 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_41
timestamp 1701704242
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1701704242
transform -1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_42
timestamp 1701704242
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1701704242
transform -1 0 23828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_43
timestamp 1701704242
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1701704242
transform -1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_44
timestamp 1701704242
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1701704242
transform -1 0 23828 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_45
timestamp 1701704242
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1701704242
transform -1 0 23828 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_46
timestamp 1701704242
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1701704242
transform -1 0 23828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_47
timestamp 1701704242
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1701704242
transform -1 0 23828 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_48
timestamp 1701704242
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1701704242
transform -1 0 23828 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_49
timestamp 1701704242
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1701704242
transform -1 0 23828 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_50
timestamp 1701704242
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1701704242
transform -1 0 23828 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_51
timestamp 1701704242
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1701704242
transform -1 0 23828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_52
timestamp 1701704242
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1701704242
transform -1 0 23828 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_53
timestamp 1701704242
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1701704242
transform -1 0 23828 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_54
timestamp 1701704242
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1701704242
transform -1 0 23828 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_55
timestamp 1701704242
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1701704242
transform -1 0 23828 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_56
timestamp 1701704242
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1701704242
transform -1 0 23828 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_57
timestamp 1701704242
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1701704242
transform -1 0 23828 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_58
timestamp 1701704242
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1701704242
transform -1 0 23828 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_59
timestamp 1701704242
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1701704242
transform -1 0 23828 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_60
timestamp 1701704242
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1701704242
transform -1 0 23828 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_61
timestamp 1701704242
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1701704242
transform -1 0 23828 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_62
timestamp 1701704242
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1701704242
transform -1 0 23828 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_63
timestamp 1701704242
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1701704242
transform -1 0 23828 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_64
timestamp 1701704242
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1701704242
transform -1 0 23828 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_65
timestamp 1701704242
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1701704242
transform -1 0 23828 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_66
timestamp 1701704242
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1701704242
transform -1 0 23828 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_67
timestamp 1701704242
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1701704242
transform -1 0 23828 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_68
timestamp 1701704242
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1701704242
transform -1 0 23828 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_69
timestamp 1701704242
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1701704242
transform -1 0 23828 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_70
timestamp 1701704242
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1701704242
transform -1 0 23828 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_71
timestamp 1701704242
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1701704242
transform -1 0 23828 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_72
timestamp 1701704242
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1701704242
transform -1 0 23828 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_73
timestamp 1701704242
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1701704242
transform -1 0 23828 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_74
timestamp 1701704242
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1701704242
transform -1 0 23828 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_75
timestamp 1701704242
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1701704242
transform -1 0 23828 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_76
timestamp 1701704242
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1701704242
transform -1 0 23828 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_77
timestamp 1701704242
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1701704242
transform -1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_78
timestamp 1701704242
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1701704242
transform -1 0 23828 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_79
timestamp 1701704242
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1701704242
transform -1 0 23828 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_80
timestamp 1701704242
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1701704242
transform -1 0 23828 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_81
timestamp 1701704242
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1701704242
transform -1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_82 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_83
timestamp 1701704242
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84
timestamp 1701704242
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 1701704242
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 1701704242
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 1701704242
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1701704242
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_89
timestamp 1701704242
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_90
timestamp 1701704242
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_91
timestamp 1701704242
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 1701704242
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 1701704242
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_94
timestamp 1701704242
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_95
timestamp 1701704242
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 1701704242
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 1701704242
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_98
timestamp 1701704242
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_99
timestamp 1701704242
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 1701704242
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 1701704242
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_102
timestamp 1701704242
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_103
timestamp 1701704242
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_104
timestamp 1701704242
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 1701704242
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_106
timestamp 1701704242
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_107
timestamp 1701704242
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_108
timestamp 1701704242
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_109
timestamp 1701704242
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_110
timestamp 1701704242
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_111
timestamp 1701704242
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_112
timestamp 1701704242
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_113
timestamp 1701704242
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_114
timestamp 1701704242
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_115
timestamp 1701704242
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 1701704242
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_117
timestamp 1701704242
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_118
timestamp 1701704242
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_119
timestamp 1701704242
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 1701704242
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 1701704242
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_122
timestamp 1701704242
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_123
timestamp 1701704242
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 1701704242
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 1701704242
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_126
timestamp 1701704242
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_127
timestamp 1701704242
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 1701704242
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 1701704242
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_130
timestamp 1701704242
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_131
timestamp 1701704242
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_132
timestamp 1701704242
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_133
timestamp 1701704242
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_134
timestamp 1701704242
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_135
timestamp 1701704242
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_136
timestamp 1701704242
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_137
timestamp 1701704242
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_138
timestamp 1701704242
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_139
timestamp 1701704242
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_140
timestamp 1701704242
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_141
timestamp 1701704242
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_142
timestamp 1701704242
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_143
timestamp 1701704242
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_144
timestamp 1701704242
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_145
timestamp 1701704242
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_146
timestamp 1701704242
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_147
timestamp 1701704242
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_148
timestamp 1701704242
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_149
timestamp 1701704242
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_150
timestamp 1701704242
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_151
timestamp 1701704242
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_152
timestamp 1701704242
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_153
timestamp 1701704242
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_154
timestamp 1701704242
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_155
timestamp 1701704242
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_156
timestamp 1701704242
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_157
timestamp 1701704242
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_158
timestamp 1701704242
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_159
timestamp 1701704242
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_160
timestamp 1701704242
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_161
timestamp 1701704242
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_162
timestamp 1701704242
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_163
timestamp 1701704242
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_164
timestamp 1701704242
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_165
timestamp 1701704242
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_166
timestamp 1701704242
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_167
timestamp 1701704242
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_168
timestamp 1701704242
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_169
timestamp 1701704242
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_170
timestamp 1701704242
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_171
timestamp 1701704242
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_172
timestamp 1701704242
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_173
timestamp 1701704242
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_174
timestamp 1701704242
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_175
timestamp 1701704242
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_176
timestamp 1701704242
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_177
timestamp 1701704242
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_178
timestamp 1701704242
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_179
timestamp 1701704242
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_180
timestamp 1701704242
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_181
timestamp 1701704242
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_182
timestamp 1701704242
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_183
timestamp 1701704242
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_184
timestamp 1701704242
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_185
timestamp 1701704242
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_186
timestamp 1701704242
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_187
timestamp 1701704242
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_188
timestamp 1701704242
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_189
timestamp 1701704242
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_190
timestamp 1701704242
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_191
timestamp 1701704242
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_192
timestamp 1701704242
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_193
timestamp 1701704242
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_194
timestamp 1701704242
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_195
timestamp 1701704242
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_196
timestamp 1701704242
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_197
timestamp 1701704242
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_198
timestamp 1701704242
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_199
timestamp 1701704242
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_200
timestamp 1701704242
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_201
timestamp 1701704242
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_202
timestamp 1701704242
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_203
timestamp 1701704242
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_204
timestamp 1701704242
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_205
timestamp 1701704242
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_206
timestamp 1701704242
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_207
timestamp 1701704242
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_208
timestamp 1701704242
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_209
timestamp 1701704242
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_210
timestamp 1701704242
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_211
timestamp 1701704242
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_212
timestamp 1701704242
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_213
timestamp 1701704242
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_214
timestamp 1701704242
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_215
timestamp 1701704242
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_216
timestamp 1701704242
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_217
timestamp 1701704242
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_218
timestamp 1701704242
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_219
timestamp 1701704242
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_220
timestamp 1701704242
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_221
timestamp 1701704242
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_222
timestamp 1701704242
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_223
timestamp 1701704242
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_224
timestamp 1701704242
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_225
timestamp 1701704242
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_226
timestamp 1701704242
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_227
timestamp 1701704242
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_228
timestamp 1701704242
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_229
timestamp 1701704242
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_230
timestamp 1701704242
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_231
timestamp 1701704242
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_232
timestamp 1701704242
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_233
timestamp 1701704242
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_234
timestamp 1701704242
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_235
timestamp 1701704242
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_236
timestamp 1701704242
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_237
timestamp 1701704242
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_238
timestamp 1701704242
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_239
timestamp 1701704242
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_240
timestamp 1701704242
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_241
timestamp 1701704242
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_242
timestamp 1701704242
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_243
timestamp 1701704242
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_244
timestamp 1701704242
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_245
timestamp 1701704242
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_246
timestamp 1701704242
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_247
timestamp 1701704242
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_248
timestamp 1701704242
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_249
timestamp 1701704242
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_250
timestamp 1701704242
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_251
timestamp 1701704242
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_252
timestamp 1701704242
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_253
timestamp 1701704242
transform 1 0 21712 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 MEM_WRITE[0]
port 0 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 MEM_WRITE[10]
port 1 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 MEM_WRITE[11]
port 2 nsew signal tristate
flabel metal2 s 10966 26344 11022 27144 0 FreeSans 224 90 0 0 MEM_WRITE[12]
port 3 nsew signal tristate
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 MEM_WRITE[13]
port 4 nsew signal tristate
flabel metal2 s 8390 26344 8446 27144 0 FreeSans 224 90 0 0 MEM_WRITE[14]
port 5 nsew signal tristate
flabel metal2 s 7746 26344 7802 27144 0 FreeSans 224 90 0 0 MEM_WRITE[15]
port 6 nsew signal tristate
flabel metal2 s 13542 26344 13598 27144 0 FreeSans 224 90 0 0 MEM_WRITE[16]
port 7 nsew signal tristate
flabel metal2 s 14186 26344 14242 27144 0 FreeSans 224 90 0 0 MEM_WRITE[17]
port 8 nsew signal tristate
flabel metal3 s 24200 13608 25000 13728 0 FreeSans 480 0 0 0 MEM_WRITE[18]
port 9 nsew signal tristate
flabel metal2 s 14830 26344 14886 27144 0 FreeSans 224 90 0 0 MEM_WRITE[19]
port 10 nsew signal tristate
flabel metal3 s 24200 12248 25000 12368 0 FreeSans 480 0 0 0 MEM_WRITE[1]
port 11 nsew signal tristate
flabel metal3 s 24200 19048 25000 19168 0 FreeSans 480 0 0 0 MEM_WRITE[20]
port 12 nsew signal tristate
flabel metal3 s 24200 18368 25000 18488 0 FreeSans 480 0 0 0 MEM_WRITE[21]
port 13 nsew signal tristate
flabel metal3 s 24200 16328 25000 16448 0 FreeSans 480 0 0 0 MEM_WRITE[22]
port 14 nsew signal tristate
flabel metal3 s 24200 15648 25000 15768 0 FreeSans 480 0 0 0 MEM_WRITE[23]
port 15 nsew signal tristate
flabel metal3 s 24200 12928 25000 13048 0 FreeSans 480 0 0 0 MEM_WRITE[24]
port 16 nsew signal tristate
flabel metal3 s 24200 14288 25000 14408 0 FreeSans 480 0 0 0 MEM_WRITE[25]
port 17 nsew signal tristate
flabel metal3 s 24200 10888 25000 11008 0 FreeSans 480 0 0 0 MEM_WRITE[26]
port 18 nsew signal tristate
flabel metal3 s 24200 11568 25000 11688 0 FreeSans 480 0 0 0 MEM_WRITE[27]
port 19 nsew signal tristate
flabel metal3 s 24200 8848 25000 8968 0 FreeSans 480 0 0 0 MEM_WRITE[28]
port 20 nsew signal tristate
flabel metal3 s 24200 8168 25000 8288 0 FreeSans 480 0 0 0 MEM_WRITE[29]
port 21 nsew signal tristate
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 MEM_WRITE[2]
port 22 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 MEM_WRITE[30]
port 23 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 MEM_WRITE[31]
port 24 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 MEM_WRITE[3]
port 25 nsew signal tristate
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 MEM_WRITE[4]
port 26 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 MEM_WRITE[5]
port 27 nsew signal tristate
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 MEM_WRITE[6]
port 28 nsew signal tristate
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 MEM_WRITE[7]
port 29 nsew signal tristate
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 MEM_WRITE[8]
port 30 nsew signal tristate
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 MEM_WRITE[9]
port 31 nsew signal tristate
flabel metal4 s -1076 -4 -756 26660 0 FreeSans 1920 90 0 0 VGND
port 32 nsew ground bidirectional
flabel metal5 s -1076 -4 26008 316 0 FreeSans 2560 0 0 0 VGND
port 32 nsew ground bidirectional
flabel metal5 s -1076 26340 26008 26660 0 FreeSans 2560 0 0 0 VGND
port 32 nsew ground bidirectional
flabel metal4 s 25688 -4 26008 26660 0 FreeSans 1920 90 0 0 VGND
port 32 nsew ground bidirectional
flabel metal4 s 2644 -4 3044 26660 0 FreeSans 1920 90 0 0 VGND
port 32 nsew ground bidirectional
flabel metal4 s 8644 -4 9044 26660 0 FreeSans 1920 90 0 0 VGND
port 32 nsew ground bidirectional
flabel metal4 s 14644 -4 15044 26660 0 FreeSans 1920 90 0 0 VGND
port 32 nsew ground bidirectional
flabel metal4 s 20644 -4 21044 26660 0 FreeSans 1920 90 0 0 VGND
port 32 nsew ground bidirectional
flabel metal5 s -1076 3716 26008 4116 0 FreeSans 2560 0 0 0 VGND
port 32 nsew ground bidirectional
flabel metal5 s -1076 9716 26008 10116 0 FreeSans 2560 0 0 0 VGND
port 32 nsew ground bidirectional
flabel metal5 s -1076 15716 26008 16116 0 FreeSans 2560 0 0 0 VGND
port 32 nsew ground bidirectional
flabel metal5 s -1076 21716 26008 22116 0 FreeSans 2560 0 0 0 VGND
port 32 nsew ground bidirectional
flabel metal4 s -416 656 -96 26000 0 FreeSans 1920 90 0 0 VPWR
port 33 nsew power bidirectional
flabel metal5 s -416 656 25348 976 0 FreeSans 2560 0 0 0 VPWR
port 33 nsew power bidirectional
flabel metal5 s -416 25680 25348 26000 0 FreeSans 2560 0 0 0 VPWR
port 33 nsew power bidirectional
flabel metal4 s 25028 656 25348 26000 0 FreeSans 1920 90 0 0 VPWR
port 33 nsew power bidirectional
flabel metal4 s 1904 -4 2304 26660 0 FreeSans 1920 90 0 0 VPWR
port 33 nsew power bidirectional
flabel metal4 s 7904 -4 8304 26660 0 FreeSans 1920 90 0 0 VPWR
port 33 nsew power bidirectional
flabel metal4 s 13904 -4 14304 26660 0 FreeSans 1920 90 0 0 VPWR
port 33 nsew power bidirectional
flabel metal4 s 19904 -4 20304 26660 0 FreeSans 1920 90 0 0 VPWR
port 33 nsew power bidirectional
flabel metal5 s -1076 2976 26008 3376 0 FreeSans 2560 0 0 0 VPWR
port 33 nsew power bidirectional
flabel metal5 s -1076 8976 26008 9376 0 FreeSans 2560 0 0 0 VPWR
port 33 nsew power bidirectional
flabel metal5 s -1076 14976 26008 15376 0 FreeSans 2560 0 0 0 VPWR
port 33 nsew power bidirectional
flabel metal5 s -1076 20976 26008 21376 0 FreeSans 2560 0 0 0 VPWR
port 33 nsew power bidirectional
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 clk
port 34 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 rst
port 35 nsew signal input
rlabel metal1 12466 23936 12466 23936 0 VGND
rlabel metal1 12466 24480 12466 24480 0 VPWR
rlabel metal1 13202 7378 13202 7378 0 ALUData1Mux.in1\[0\]
rlabel metal1 6036 18258 6036 18258 0 ALUData1Mux.in1\[10\]
rlabel metal1 2553 14450 2553 14450 0 ALUData1Mux.in1\[11\]
rlabel metal1 7452 15674 7452 15674 0 ALUData1Mux.in1\[12\]
rlabel metal1 11362 12172 11362 12172 0 ALUData1Mux.in1\[13\]
rlabel metal1 6936 20910 6936 20910 0 ALUData1Mux.in1\[14\]
rlabel metal1 5520 20026 5520 20026 0 ALUData1Mux.in1\[15\]
rlabel metal1 12732 21522 12732 21522 0 ALUData1Mux.in1\[16\]
rlabel via1 11817 20502 11817 20502 0 ALUData1Mux.in1\[17\]
rlabel metal1 13432 14042 13432 14042 0 ALUData1Mux.in1\[18\]
rlabel metal2 13294 17748 13294 17748 0 ALUData1Mux.in1\[19\]
rlabel metal1 13160 11118 13160 11118 0 ALUData1Mux.in1\[1\]
rlabel metal1 18528 19346 18528 19346 0 ALUData1Mux.in1\[20\]
rlabel metal1 17935 20502 17935 20502 0 ALUData1Mux.in1\[21\]
rlabel metal1 20060 16490 20060 16490 0 ALUData1Mux.in1\[22\]
rlabel metal2 17066 15096 17066 15096 0 ALUData1Mux.in1\[23\]
rlabel metal1 22172 13498 22172 13498 0 ALUData1Mux.in1\[24\]
rlabel metal1 20930 14518 20930 14518 0 ALUData1Mux.in1\[25\]
rlabel metal1 21850 8262 21850 8262 0 ALUData1Mux.in1\[26\]
rlabel metal1 17710 9010 17710 9010 0 ALUData1Mux.in1\[27\]
rlabel metal1 19872 8262 19872 8262 0 ALUData1Mux.in1\[28\]
rlabel via1 21482 7242 21482 7242 0 ALUData1Mux.in1\[29\]
rlabel metal1 10350 4998 10350 4998 0 ALUData1Mux.in1\[2\]
rlabel metal1 17081 6698 17081 6698 0 ALUData1Mux.in1\[30\]
rlabel metal1 18216 5134 18216 5134 0 ALUData1Mux.in1\[31\]
rlabel via1 12654 4182 12654 4182 0 ALUData1Mux.in1\[3\]
rlabel via1 4630 5610 4630 5610 0 ALUData1Mux.in1\[4\]
rlabel metal1 3721 6290 3721 6290 0 ALUData1Mux.in1\[5\]
rlabel metal2 2990 9214 2990 9214 0 ALUData1Mux.in1\[6\]
rlabel metal1 10258 9146 10258 9146 0 ALUData1Mux.in1\[7\]
rlabel metal1 5004 12818 5004 12818 0 ALUData1Mux.in1\[8\]
rlabel metal1 1610 10132 1610 10132 0 ALUData1Mux.in1\[9\]
rlabel metal2 12558 9316 12558 9316 0 ALUData1Mux.in2\[0\]
rlabel metal1 3358 15470 3358 15470 0 ALUData1Mux.in2\[10\]
rlabel metal1 7452 15130 7452 15130 0 ALUData1Mux.in2\[11\]
rlabel metal1 11270 17850 11270 17850 0 ALUData1Mux.in2\[12\]
rlabel metal2 11362 15402 11362 15402 0 ALUData1Mux.in2\[13\]
rlabel metal1 10166 20570 10166 20570 0 ALUData1Mux.in2\[14\]
rlabel metal1 9660 19142 9660 19142 0 ALUData1Mux.in2\[15\]
rlabel metal1 17296 20978 17296 20978 0 ALUData1Mux.in2\[16\]
rlabel metal1 16560 20570 16560 20570 0 ALUData1Mux.in2\[17\]
rlabel metal1 12328 14994 12328 14994 0 ALUData1Mux.in2\[18\]
rlabel metal1 12282 16660 12282 16660 0 ALUData1Mux.in2\[19\]
rlabel metal1 12282 10540 12282 10540 0 ALUData1Mux.in2\[1\]
rlabel metal1 17526 18734 17526 18734 0 ALUData1Mux.in2\[20\]
rlabel metal1 16054 19210 16054 19210 0 ALUData1Mux.in2\[21\]
rlabel metal1 19182 13838 19182 13838 0 ALUData1Mux.in2\[22\]
rlabel metal1 19688 14790 19688 14790 0 ALUData1Mux.in2\[23\]
rlabel metal1 21298 10574 21298 10574 0 ALUData1Mux.in2\[24\]
rlabel metal1 21344 13838 21344 13838 0 ALUData1Mux.in2\[25\]
rlabel metal2 21850 6834 21850 6834 0 ALUData1Mux.in2\[26\]
rlabel metal1 16974 8466 16974 8466 0 ALUData1Mux.in2\[27\]
rlabel metal1 20930 5814 20930 5814 0 ALUData1Mux.in2\[28\]
rlabel metal1 21160 6290 21160 6290 0 ALUData1Mux.in2\[29\]
rlabel metal1 9936 3502 9936 3502 0 ALUData1Mux.in2\[2\]
rlabel metal2 16146 7004 16146 7004 0 ALUData1Mux.in2\[30\]
rlabel metal1 14536 7514 14536 7514 0 ALUData1Mux.in2\[31\]
rlabel metal1 7176 4046 7176 4046 0 ALUData1Mux.in2\[3\]
rlabel metal1 9154 4046 9154 4046 0 ALUData1Mux.in2\[4\]
rlabel metal1 9660 6086 9660 6086 0 ALUData1Mux.in2\[5\]
rlabel metal1 7728 8466 7728 8466 0 ALUData1Mux.in2\[6\]
rlabel metal1 11224 6290 11224 6290 0 ALUData1Mux.in2\[7\]
rlabel metal1 8648 10574 8648 10574 0 ALUData1Mux.in2\[8\]
rlabel metal1 7130 12818 7130 12818 0 ALUData1Mux.in2\[9\]
rlabel metal2 13570 8194 13570 8194 0 ALUData1Mux.in3\[0\]
rlabel metal1 3220 16082 3220 16082 0 ALUData1Mux.in3\[10\]
rlabel metal1 4232 14382 4232 14382 0 ALUData1Mux.in3\[11\]
rlabel metal1 6578 15878 6578 15878 0 ALUData1Mux.in3\[12\]
rlabel metal1 11316 13294 11316 13294 0 ALUData1Mux.in3\[13\]
rlabel metal1 8142 20026 8142 20026 0 ALUData1Mux.in3\[14\]
rlabel metal1 7360 20230 7360 20230 0 ALUData1Mux.in3\[15\]
rlabel metal1 15548 21114 15548 21114 0 ALUData1Mux.in3\[16\]
rlabel metal1 14444 20298 14444 20298 0 ALUData1Mux.in3\[17\]
rlabel metal1 13616 15674 13616 15674 0 ALUData1Mux.in3\[18\]
rlabel metal1 13432 17850 13432 17850 0 ALUData1Mux.in3\[19\]
rlabel metal1 13800 10234 13800 10234 0 ALUData1Mux.in3\[1\]
rlabel metal1 21160 18394 21160 18394 0 ALUData1Mux.in3\[20\]
rlabel metal1 20562 18938 20562 18938 0 ALUData1Mux.in3\[21\]
rlabel metal1 21551 14858 21551 14858 0 ALUData1Mux.in3\[22\]
rlabel metal1 16192 13906 16192 13906 0 ALUData1Mux.in3\[23\]
rlabel metal2 23000 14348 23000 14348 0 ALUData1Mux.in3\[24\]
rlabel metal2 22126 15572 22126 15572 0 ALUData1Mux.in3\[25\]
rlabel metal1 22218 4658 22218 4658 0 ALUData1Mux.in3\[26\]
rlabel metal1 17710 12954 17710 12954 0 ALUData1Mux.in3\[27\]
rlabel metal2 22586 5372 22586 5372 0 ALUData1Mux.in3\[28\]
rlabel metal2 23506 5916 23506 5916 0 ALUData1Mux.in3\[29\]
rlabel metal1 9517 5270 9517 5270 0 ALUData1Mux.in3\[2\]
rlabel metal1 19826 7990 19826 7990 0 ALUData1Mux.in3\[30\]
rlabel metal1 17112 5202 17112 5202 0 ALUData1Mux.in3\[31\]
rlabel metal1 12052 5066 12052 5066 0 ALUData1Mux.in3\[3\]
rlabel metal1 7866 4590 7866 4590 0 ALUData1Mux.in3\[4\]
rlabel metal2 6670 5338 6670 5338 0 ALUData1Mux.in3\[5\]
rlabel metal1 2346 8296 2346 8296 0 ALUData1Mux.in3\[6\]
rlabel metal1 2438 7820 2438 7820 0 ALUData1Mux.in3\[7\]
rlabel metal1 3726 10030 3726 10030 0 ALUData1Mux.in3\[8\]
rlabel metal1 2438 11084 2438 11084 0 ALUData1Mux.in3\[9\]
rlabel metal2 12098 7548 12098 7548 0 EX_MEM.i_ALUresult\[0\]
rlabel metal1 4998 16150 4998 16150 0 EX_MEM.i_ALUresult\[10\]
rlabel via1 6490 14382 6490 14382 0 EX_MEM.i_ALUresult\[11\]
rlabel via1 7870 16082 7870 16082 0 EX_MEM.i_ALUresult\[12\]
rlabel metal3 9614 12580 9614 12580 0 EX_MEM.i_ALUresult\[13\]
rlabel metal1 8008 19754 8008 19754 0 EX_MEM.i_ALUresult\[14\]
rlabel metal1 7962 20434 7962 20434 0 EX_MEM.i_ALUresult\[15\]
rlabel metal1 14066 20910 14066 20910 0 EX_MEM.i_ALUresult\[16\]
rlabel metal1 13192 20434 13192 20434 0 EX_MEM.i_ALUresult\[17\]
rlabel via1 12369 15402 12369 15402 0 EX_MEM.i_ALUresult\[18\]
rlabel metal2 12098 16898 12098 16898 0 EX_MEM.i_ALUresult\[19\]
rlabel via1 12829 10030 12829 10030 0 EX_MEM.i_ALUresult\[1\]
rlabel metal1 19810 18326 19810 18326 0 EX_MEM.i_ALUresult\[20\]
rlabel metal1 19683 18666 19683 18666 0 EX_MEM.i_ALUresult\[21\]
rlabel metal1 19810 15062 19810 15062 0 EX_MEM.i_ALUresult\[22\]
rlabel metal1 15630 14382 15630 14382 0 EX_MEM.i_ALUresult\[23\]
rlabel metal1 22908 12614 22908 12614 0 EX_MEM.i_ALUresult\[24\]
rlabel metal1 23230 13872 23230 13872 0 EX_MEM.i_ALUresult\[25\]
rlabel metal1 20684 8874 20684 8874 0 EX_MEM.i_ALUresult\[26\]
rlabel metal1 19560 12818 19560 12818 0 EX_MEM.i_ALUresult\[27\]
rlabel metal1 21942 6766 21942 6766 0 EX_MEM.i_ALUresult\[28\]
rlabel metal1 23056 7378 23056 7378 0 EX_MEM.i_ALUresult\[29\]
rlabel metal1 12953 5610 12953 5610 0 EX_MEM.i_ALUresult\[2\]
rlabel metal1 15686 6630 15686 6630 0 EX_MEM.i_ALUresult\[30\]
rlabel metal1 17996 7378 17996 7378 0 EX_MEM.i_ALUresult\[31\]
rlabel metal2 12926 4556 12926 4556 0 EX_MEM.i_ALUresult\[3\]
rlabel metal1 6562 5270 6562 5270 0 EX_MEM.i_ALUresult\[4\]
rlabel metal1 4958 6290 4958 6290 0 EX_MEM.i_ALUresult\[5\]
rlabel metal1 4922 7242 4922 7242 0 EX_MEM.i_ALUresult\[6\]
rlabel metal2 8970 8228 8970 8228 0 EX_MEM.i_ALUresult\[7\]
rlabel metal2 6210 12517 6210 12517 0 EX_MEM.i_ALUresult\[8\]
rlabel metal1 4692 12614 4692 12614 0 EX_MEM.i_ALUresult\[9\]
rlabel via1 11081 5678 11081 5678 0 ID_EX.i_ReadData1_in\[0\]
rlabel metal1 5004 14994 5004 14994 0 ID_EX.i_ReadData1_in\[10\]
rlabel metal1 4738 13804 4738 13804 0 ID_EX.i_ReadData1_in\[11\]
rlabel metal1 8468 15402 8468 15402 0 ID_EX.i_ReadData1_in\[12\]
rlabel metal2 9292 13260 9292 13260 0 ID_EX.i_ReadData1_in\[13\]
rlabel metal1 5791 18734 5791 18734 0 ID_EX.i_ReadData1_in\[14\]
rlabel metal1 6444 19754 6444 19754 0 ID_EX.i_ReadData1_in\[15\]
rlabel metal2 12098 20808 12098 20808 0 ID_EX.i_ReadData1_in\[16\]
rlabel metal2 11362 20706 11362 20706 0 ID_EX.i_ReadData1_in\[17\]
rlabel metal1 12272 13906 12272 13906 0 ID_EX.i_ReadData1_in\[18\]
rlabel metal2 13202 17918 13202 17918 0 ID_EX.i_ReadData1_in\[19\]
rlabel metal1 10258 11322 10258 11322 0 ID_EX.i_ReadData1_in\[1\]
rlabel metal2 18170 18870 18170 18870 0 ID_EX.i_ReadData1_in\[20\]
rlabel metal2 18078 19074 18078 19074 0 ID_EX.i_ReadData1_in\[21\]
rlabel metal1 18680 13974 18680 13974 0 ID_EX.i_ReadData1_in\[22\]
rlabel metal1 17668 14382 17668 14382 0 ID_EX.i_ReadData1_in\[23\]
rlabel metal1 18538 12682 18538 12682 0 ID_EX.i_ReadData1_in\[24\]
rlabel metal2 19826 13634 19826 13634 0 ID_EX.i_ReadData1_in\[25\]
rlabel metal1 21206 10234 21206 10234 0 ID_EX.i_ReadData1_in\[26\]
rlabel metal1 15548 10778 15548 10778 0 ID_EX.i_ReadData1_in\[27\]
rlabel metal1 20750 8534 20750 8534 0 ID_EX.i_ReadData1_in\[28\]
rlabel metal1 19182 6630 19182 6630 0 ID_EX.i_ReadData1_in\[29\]
rlabel metal2 8418 7072 8418 7072 0 ID_EX.i_ReadData1_in\[2\]
rlabel metal1 15916 6970 15916 6970 0 ID_EX.i_ReadData1_in\[30\]
rlabel metal1 15405 5610 15405 5610 0 ID_EX.i_ReadData1_in\[31\]
rlabel metal2 9614 4505 9614 4505 0 ID_EX.i_ReadData1_in\[3\]
rlabel metal1 4544 5202 4544 5202 0 ID_EX.i_ReadData1_in\[4\]
rlabel via1 3629 8534 3629 8534 0 ID_EX.i_ReadData1_in\[5\]
rlabel metal1 3312 9350 3312 9350 0 ID_EX.i_ReadData1_in\[6\]
rlabel metal2 9890 8194 9890 8194 0 ID_EX.i_ReadData1_in\[7\]
rlabel metal1 1840 12614 1840 12614 0 ID_EX.i_ReadData1_in\[8\]
rlabel metal1 2507 13158 2507 13158 0 ID_EX.i_ReadData1_in\[9\]
rlabel metal2 12282 959 12282 959 0 MEM_WRITE[0]
rlabel metal3 820 17068 820 17068 0 MEM_WRITE[10]
rlabel metal3 820 15708 820 15708 0 MEM_WRITE[11]
rlabel metal1 11454 24242 11454 24242 0 MEM_WRITE[12]
rlabel metal3 820 13668 820 13668 0 MEM_WRITE[13]
rlabel metal1 8878 24242 8878 24242 0 MEM_WRITE[14]
rlabel metal1 7912 24242 7912 24242 0 MEM_WRITE[15]
rlabel metal1 13938 24242 13938 24242 0 MEM_WRITE[16]
rlabel metal1 14858 24174 14858 24174 0 MEM_WRITE[17]
rlabel metal2 23414 13515 23414 13515 0 MEM_WRITE[18]
rlabel metal1 15226 24242 15226 24242 0 MEM_WRITE[19]
rlabel metal1 22908 9010 22908 9010 0 MEM_WRITE[1]
rlabel metal2 23322 19227 23322 19227 0 MEM_WRITE[20]
rlabel metal2 23322 18547 23322 18547 0 MEM_WRITE[21]
rlabel metal2 23322 16745 23322 16745 0 MEM_WRITE[22]
rlabel metal1 23276 16490 23276 16490 0 MEM_WRITE[23]
rlabel metal1 22954 13226 22954 13226 0 MEM_WRITE[24]
rlabel metal1 23368 14314 23368 14314 0 MEM_WRITE[25]
rlabel metal2 22494 10489 22494 10489 0 MEM_WRITE[26]
rlabel metal2 23322 10455 23322 10455 0 MEM_WRITE[27]
rlabel metal1 23046 6834 23046 6834 0 MEM_WRITE[28]
rlabel metal2 23322 6273 23322 6273 0 MEM_WRITE[29]
rlabel metal2 13570 1554 13570 1554 0 MEM_WRITE[2]
rlabel metal2 17434 959 17434 959 0 MEM_WRITE[30]
rlabel metal2 18078 1554 18078 1554 0 MEM_WRITE[31]
rlabel metal2 12926 1554 12926 1554 0 MEM_WRITE[3]
rlabel metal2 7130 1639 7130 1639 0 MEM_WRITE[4]
rlabel metal2 7774 1554 7774 1554 0 MEM_WRITE[5]
rlabel metal3 1027 10948 1027 10948 0 MEM_WRITE[6]
rlabel metal1 11454 2958 11454 2958 0 MEM_WRITE[7]
rlabel metal3 820 12308 820 12308 0 MEM_WRITE[8]
rlabel metal3 820 12988 820 12988 0 MEM_WRITE[9]
rlabel metal2 11546 5474 11546 5474 0 _160_
rlabel metal1 10488 7990 10488 7990 0 _161_
rlabel metal1 8924 3910 8924 3910 0 _162_
rlabel metal2 7314 4573 7314 4573 0 _163_
rlabel metal1 1518 5542 1518 5542 0 _164_
rlabel metal1 3450 5338 3450 5338 0 _165_
rlabel metal2 2806 5763 2806 5763 0 _166_
rlabel metal1 5740 7854 5740 7854 0 _167_
rlabel metal2 1840 10540 1840 10540 0 _168_
rlabel metal1 3496 5542 3496 5542 0 _169_
rlabel metal2 3082 16014 3082 16014 0 _170_
rlabel via1 2157 13906 2157 13906 0 _171_
rlabel metal1 6220 16558 6220 16558 0 _172_
rlabel via1 5101 13906 5101 13906 0 _173_
rlabel metal1 4365 18734 4365 18734 0 _174_
rlabel metal1 4830 18122 4830 18122 0 _175_
rlabel metal1 12190 21896 12190 21896 0 _176_
rlabel metal1 11040 22406 11040 22406 0 _177_
rlabel via1 11090 13906 11090 13906 0 _178_
rlabel via1 10897 15470 10897 15470 0 _179_
rlabel via1 15313 17170 15313 17170 0 _180_
rlabel metal1 14704 17578 14704 17578 0 _181_
rlabel metal1 16882 14008 16882 14008 0 _182_
rlabel metal1 16422 12750 16422 12750 0 _183_
rlabel metal1 20623 13226 20623 13226 0 _184_
rlabel metal1 18032 13158 18032 13158 0 _185_
rlabel metal1 21298 9894 21298 9894 0 _186_
rlabel metal1 19320 10778 19320 10778 0 _187_
rlabel metal2 18538 7106 18538 7106 0 _188_
rlabel metal1 18906 5066 18906 5066 0 _189_
rlabel metal1 15226 5338 15226 5338 0 _190_
rlabel metal1 14076 4794 14076 4794 0 _191_
rlabel metal1 18584 14450 18584 14450 0 _192_
rlabel metal1 14490 4624 14490 4624 0 _193_
rlabel metal1 13938 5814 13938 5814 0 _194_
rlabel metal1 18216 5202 18216 5202 0 _195_
rlabel metal1 18768 6290 18768 6290 0 _196_
rlabel metal1 18400 9894 18400 9894 0 _197_
rlabel metal2 19734 11696 19734 11696 0 _198_
rlabel metal2 18998 13333 18998 13333 0 _199_
rlabel metal2 14398 13005 14398 13005 0 _200_
rlabel metal1 17020 12614 17020 12614 0 _201_
rlabel metal1 16698 13872 16698 13872 0 _202_
rlabel metal1 15962 19278 15962 19278 0 _203_
rlabel metal1 15870 19482 15870 19482 0 _204_
rlabel metal2 14628 19380 14628 19380 0 _205_
rlabel metal1 10442 17646 10442 17646 0 _206_
rlabel metal2 16330 14756 16330 14756 0 _207_
rlabel metal2 16514 21420 16514 21420 0 _208_
rlabel metal1 13892 19278 13892 19278 0 _209_
rlabel metal1 5060 18258 5060 18258 0 _210_
rlabel metal1 10810 18394 10810 18394 0 _211_
rlabel metal1 9660 14450 9660 14450 0 _212_
rlabel metal2 11546 16626 11546 16626 0 _213_
rlabel metal1 11960 12138 11960 12138 0 _214_
rlabel metal2 2254 15521 2254 15521 0 _215_
rlabel metal1 8832 16422 8832 16422 0 _216_
rlabel metal1 3174 5678 3174 5678 0 _217_
rlabel metal1 7038 9486 7038 9486 0 _218_
rlabel metal1 6026 7174 6026 7174 0 _219_
rlabel metal2 2162 5729 2162 5729 0 _220_
rlabel metal1 8740 9894 8740 9894 0 _221_
rlabel metal1 1610 5644 1610 5644 0 _222_
rlabel metal2 9062 3978 9062 3978 0 _223_
rlabel metal1 10074 4114 10074 4114 0 _224_
rlabel metal1 11684 11186 11684 11186 0 _225_
rlabel metal1 11960 7514 11960 7514 0 _226_
rlabel metal1 14812 14042 14812 14042 0 _227_
rlabel metal1 11454 10506 11454 10506 0 _228_
rlabel metal1 4600 8058 4600 8058 0 _229_
rlabel metal1 10396 17238 10396 17238 0 _230_
rlabel metal1 14674 11322 14674 11322 0 _231_
rlabel metal1 13846 5882 13846 5882 0 _232_
rlabel metal2 6854 14960 6854 14960 0 _233_
rlabel metal1 15134 15334 15134 15334 0 _234_
rlabel via2 2438 9435 2438 9435 0 _235_
rlabel metal1 10442 4794 10442 4794 0 _236_
rlabel metal1 15364 12954 15364 12954 0 _237_
rlabel metal2 16698 10166 16698 10166 0 _238_
rlabel metal2 2530 13838 2530 13838 0 _239_
rlabel metal1 14260 18258 14260 18258 0 _240_
rlabel metal1 14858 13430 14858 13430 0 _241_
rlabel metal1 9108 5882 9108 5882 0 _242_
rlabel metal1 9890 17850 9890 17850 0 _243_
rlabel metal1 14950 13158 14950 13158 0 _244_
rlabel metal2 3818 16592 3818 16592 0 clk
rlabel metal2 13570 14110 13570 14110 0 clknet_0__227_
rlabel metal1 12972 11798 12972 11798 0 clknet_0__228_
rlabel metal1 7912 8534 7912 8534 0 clknet_0__229_
rlabel metal1 7038 17238 7038 17238 0 clknet_0__230_
rlabel metal1 16376 13498 16376 13498 0 clknet_0__231_
rlabel metal1 9292 9350 9292 9350 0 clknet_0__232_
rlabel metal2 9522 17306 9522 17306 0 clknet_0__233_
rlabel metal1 18446 15470 18446 15470 0 clknet_0__234_
rlabel metal2 14214 8738 14214 8738 0 clknet_0__235_
rlabel metal1 8418 15130 8418 15130 0 clknet_0__236_
rlabel metal1 17526 17306 17526 17306 0 clknet_0__237_
rlabel metal2 17986 8908 17986 8908 0 clknet_0__238_
rlabel metal1 8786 13906 8786 13906 0 clknet_0__239_
rlabel metal1 14858 18394 14858 18394 0 clknet_0__240_
rlabel metal1 17756 11118 17756 11118 0 clknet_0__241_
rlabel metal1 9062 13158 9062 13158 0 clknet_0__242_
rlabel metal1 13984 18326 13984 18326 0 clknet_0__243_
rlabel metal2 20562 11934 20562 11934 0 clknet_0__244_
rlabel metal1 15962 9622 15962 9622 0 clknet_0_clk
rlabel metal2 9476 7956 9476 7956 0 clknet_1_0__leaf__227_
rlabel metal2 11592 13668 11592 13668 0 clknet_1_0__leaf__228_
rlabel metal2 2254 15980 2254 15980 0 clknet_1_0__leaf__229_
rlabel metal1 4278 20876 4278 20876 0 clknet_1_0__leaf__230_
rlabel metal1 16560 12070 16560 12070 0 clknet_1_0__leaf__231_
rlabel metal1 1794 8500 1794 8500 0 clknet_1_0__leaf__232_
rlabel metal2 12190 7905 12190 7905 0 clknet_1_0__leaf__233_
rlabel metal1 17204 15130 17204 15130 0 clknet_1_0__leaf__234_
rlabel metal1 13524 4590 13524 4590 0 clknet_1_0__leaf__235_
rlabel metal1 1748 7378 1748 7378 0 clknet_1_0__leaf__236_
rlabel metal1 16238 16116 16238 16116 0 clknet_1_0__leaf__237_
rlabel metal1 13938 10642 13938 10642 0 clknet_1_0__leaf__238_
rlabel metal1 6992 10438 6992 10438 0 clknet_1_0__leaf__239_
rlabel metal1 14398 21556 14398 21556 0 clknet_1_0__leaf__240_
rlabel metal1 14398 12886 14398 12886 0 clknet_1_0__leaf__241_
rlabel metal1 12098 3468 12098 3468 0 clknet_1_0__leaf__242_
rlabel metal1 6716 20434 6716 20434 0 clknet_1_0__leaf__243_
rlabel metal2 16744 14212 16744 14212 0 clknet_1_0__leaf__244_
rlabel metal1 14398 13328 14398 13328 0 clknet_1_1__leaf__227_
rlabel metal2 13616 12818 13616 12818 0 clknet_1_1__leaf__228_
rlabel metal2 14398 8534 14398 8534 0 clknet_1_1__leaf__229_
rlabel metal1 2277 12818 2277 12818 0 clknet_1_1__leaf__230_
rlabel metal1 18998 13260 18998 13260 0 clknet_1_1__leaf__231_
rlabel metal1 14398 7854 14398 7854 0 clknet_1_1__leaf__232_
rlabel metal1 6394 20434 6394 20434 0 clknet_1_1__leaf__233_
rlabel metal1 18814 17680 18814 17680 0 clknet_1_1__leaf__234_
rlabel metal1 15962 9554 15962 9554 0 clknet_1_1__leaf__235_
rlabel metal1 6394 19380 6394 19380 0 clknet_1_1__leaf__236_
rlabel metal1 17986 20944 17986 20944 0 clknet_1_1__leaf__237_
rlabel metal1 21574 7412 21574 7412 0 clknet_1_1__leaf__238_
rlabel metal1 1610 15062 1610 15062 0 clknet_1_1__leaf__239_
rlabel metal1 17020 17510 17020 17510 0 clknet_1_1__leaf__240_
rlabel metal1 21804 11186 21804 11186 0 clknet_1_1__leaf__241_
rlabel metal1 4370 15470 4370 15470 0 clknet_1_1__leaf__242_
rlabel metal1 14444 16082 14444 16082 0 clknet_1_1__leaf__243_
rlabel metal1 21574 16116 21574 16116 0 clknet_1_1__leaf__244_
rlabel metal1 1886 6154 1886 6154 0 clknet_3_0__leaf_clk
rlabel metal1 7038 7412 7038 7412 0 clknet_3_1__leaf_clk
rlabel metal1 6716 20978 6716 20978 0 clknet_3_2__leaf_clk
rlabel metal1 9752 14382 9752 14382 0 clknet_3_3__leaf_clk
rlabel metal1 14122 6154 14122 6154 0 clknet_3_4__leaf_clk
rlabel metal1 21804 12614 21804 12614 0 clknet_3_5__leaf_clk
rlabel metal1 13662 16082 13662 16082 0 clknet_3_6__leaf_clk
rlabel metal1 21804 13906 21804 13906 0 clknet_3_7__leaf_clk
rlabel metal1 11270 2482 11270 2482 0 net1
rlabel metal1 14628 24174 14628 24174 0 net10
rlabel metal2 3174 6460 3174 6460 0 net100
rlabel metal2 2806 6919 2806 6919 0 net101
rlabel metal1 1518 10574 1518 10574 0 net102
rlabel metal1 1564 6426 1564 6426 0 net103
rlabel metal2 1886 15164 1886 15164 0 net104
rlabel metal1 1840 13906 1840 13906 0 net105
rlabel metal1 6624 16626 6624 16626 0 net106
rlabel metal2 4830 13396 4830 13396 0 net107
rlabel metal1 4002 18394 4002 18394 0 net108
rlabel metal1 4462 20910 4462 20910 0 net109
rlabel metal1 15502 14280 15502 14280 0 net11
rlabel metal1 9522 20910 9522 20910 0 net110
rlabel metal1 11086 19890 11086 19890 0 net111
rlabel metal1 8924 12954 8924 12954 0 net112
rlabel metal1 10580 15538 10580 15538 0 net113
rlabel metal1 15042 17204 15042 17204 0 net114
rlabel metal1 15686 17646 15686 17646 0 net115
rlabel metal1 17710 15606 17710 15606 0 net116
rlabel metal1 15870 12852 15870 12852 0 net117
rlabel metal1 20010 13294 20010 13294 0 net118
rlabel metal1 17066 10778 17066 10778 0 net119
rlabel metal1 15364 24174 15364 24174 0 net12
rlabel metal1 20286 10540 20286 10540 0 net120
rlabel metal1 15594 12206 15594 12206 0 net121
rlabel metal1 18860 6970 18860 6970 0 net122
rlabel metal1 19918 9452 19918 9452 0 net123
rlabel metal1 14076 7854 14076 7854 0 net124
rlabel metal1 14398 5270 14398 5270 0 net125
rlabel metal1 10672 4114 10672 4114 0 net126
rlabel metal1 11224 12750 11224 12750 0 net127
rlabel metal1 11638 3706 11638 3706 0 net128
rlabel metal1 9890 3706 9890 3706 0 net129
rlabel metal1 21114 8840 21114 8840 0 net13
rlabel metal1 3956 5134 3956 5134 0 net130
rlabel metal1 3128 5882 3128 5882 0 net131
rlabel metal1 2300 11118 2300 11118 0 net132
rlabel metal2 9246 8772 9246 8772 0 net133
rlabel metal1 1656 6834 1656 6834 0 net134
rlabel metal2 3082 9554 3082 9554 0 net135
rlabel metal1 4508 14994 4508 14994 0 net136
rlabel metal1 3634 14450 3634 14450 0 net137
rlabel metal1 8786 15606 8786 15606 0 net138
rlabel metal1 10856 8058 10856 8058 0 net139
rlabel metal2 21390 19584 21390 19584 0 net14
rlabel metal1 4876 18394 4876 18394 0 net140
rlabel metal1 6762 19958 6762 19958 0 net141
rlabel metal1 9292 18938 9292 18938 0 net142
rlabel metal1 11086 21046 11086 21046 0 net143
rlabel metal1 13386 13430 13386 13430 0 net144
rlabel metal1 11684 17102 11684 17102 0 net145
rlabel metal1 18538 18938 18538 18938 0 net146
rlabel metal1 18630 17850 18630 17850 0 net147
rlabel metal1 19090 13940 19090 13940 0 net148
rlabel metal1 18446 14518 18446 14518 0 net149
rlabel metal2 21482 19482 21482 19482 0 net15
rlabel metal1 21160 13294 21160 13294 0 net150
rlabel metal1 20930 12614 20930 12614 0 net151
rlabel metal1 23230 10778 23230 10778 0 net152
rlabel metal2 16238 10064 16238 10064 0 net153
rlabel metal1 21206 8500 21206 8500 0 net154
rlabel metal1 19504 5882 19504 5882 0 net155
rlabel metal1 16192 5338 16192 5338 0 net156
rlabel metal2 15686 5508 15686 5508 0 net157
rlabel metal1 15962 7514 15962 7514 0 net158
rlabel metal1 14306 9486 14306 9486 0 net159
rlabel metal1 21735 17034 21735 17034 0 net16
rlabel metal2 12466 5236 12466 5236 0 net160
rlabel metal1 13156 4658 13156 4658 0 net161
rlabel metal1 4002 5882 4002 5882 0 net162
rlabel metal2 5842 5780 5842 5780 0 net163
rlabel metal1 5888 3978 5888 3978 0 net164
rlabel metal1 8740 9146 8740 9146 0 net165
rlabel metal2 2622 15708 2622 15708 0 net166
rlabel metal1 3358 7208 3358 7208 0 net167
rlabel metal1 4370 15674 4370 15674 0 net168
rlabel metal1 4370 15538 4370 15538 0 net169
rlabel metal1 18768 14790 18768 14790 0 net17
rlabel metal1 9430 19346 9430 19346 0 net170
rlabel metal1 13294 13498 13294 13498 0 net171
rlabel metal2 6854 20332 6854 20332 0 net172
rlabel metal1 6578 19346 6578 19346 0 net173
rlabel metal1 13892 19822 13892 19822 0 net174
rlabel metal2 12558 20366 12558 20366 0 net175
rlabel metal1 13616 14450 13616 14450 0 net176
rlabel metal1 13386 17204 13386 17204 0 net177
rlabel metal1 19320 19822 19320 19822 0 net178
rlabel metal1 18492 20434 18492 20434 0 net179
rlabel metal1 20608 11526 20608 11526 0 net18
rlabel metal1 20010 17204 20010 17204 0 net180
rlabel metal1 16652 14994 16652 14994 0 net181
rlabel metal1 21390 11594 21390 11594 0 net182
rlabel metal1 22770 14042 22770 14042 0 net183
rlabel metal2 21482 8772 21482 8772 0 net184
rlabel metal2 21114 11968 21114 11968 0 net185
rlabel metal1 20286 6426 20286 6426 0 net186
rlabel metal1 20378 6188 20378 6188 0 net187
rlabel metal1 18630 5338 18630 5338 0 net188
rlabel metal1 16790 4794 16790 4794 0 net189
rlabel metal1 22034 14416 22034 14416 0 net19
rlabel metal2 13110 5984 13110 5984 0 net190
rlabel metal2 12558 10234 12558 10234 0 net191
rlabel metal1 14444 5338 14444 5338 0 net192
rlabel metal1 13432 4250 13432 4250 0 net193
rlabel metal1 11730 13770 11730 13770 0 net194
rlabel metal2 15778 13328 15778 13328 0 net195
rlabel metal2 9430 4182 9430 4182 0 net196
rlabel metal1 9292 4114 9292 4114 0 net197
rlabel metal2 11914 8296 11914 8296 0 net198
rlabel metal1 11684 3502 11684 3502 0 net199
rlabel metal2 12604 6324 12604 6324 0 net2
rlabel metal1 22172 10030 22172 10030 0 net20
rlabel metal1 14582 5814 14582 5814 0 net200
rlabel metal1 14490 8364 14490 8364 0 net201
rlabel metal1 11776 15946 11776 15946 0 net202
rlabel metal2 6762 17782 6762 17782 0 net203
rlabel metal2 11638 17272 11638 17272 0 net204
rlabel metal1 10304 17510 10304 17510 0 net205
rlabel metal1 8878 3638 8878 3638 0 net206
rlabel metal1 7636 4114 7636 4114 0 net207
rlabel metal1 16560 19210 16560 19210 0 net208
rlabel metal1 14444 18734 14444 18734 0 net209
rlabel metal1 22816 10030 22816 10030 0 net21
rlabel metal1 17618 8466 17618 8466 0 net210
rlabel metal1 20884 10642 20884 10642 0 net211
rlabel metal1 10534 15946 10534 15946 0 net212
rlabel metal1 1656 10642 1656 10642 0 net213
rlabel metal1 11454 11254 11454 11254 0 net214
rlabel metal1 10718 7854 10718 7854 0 net215
rlabel metal1 14628 17782 14628 17782 0 net216
rlabel metal1 5382 16490 5382 16490 0 net217
rlabel metal1 8418 9486 8418 9486 0 net218
rlabel metal1 1426 6800 1426 6800 0 net219
rlabel metal1 22034 6698 22034 6698 0 net22
rlabel metal1 16560 20298 16560 20298 0 net220
rlabel metal2 16238 14552 16238 14552 0 net221
rlabel metal1 9982 7446 9982 7446 0 net222
rlabel metal1 3772 15674 3772 15674 0 net223
rlabel metal1 14214 19176 14214 19176 0 net224
rlabel metal1 11454 18122 11454 18122 0 net225
rlabel metal1 9338 6902 9338 6902 0 net226
rlabel metal1 19964 11254 19964 11254 0 net227
rlabel metal1 8970 8330 8970 8330 0 net228
rlabel metal1 17802 8296 17802 8296 0 net229
rlabel metal1 21022 5746 21022 5746 0 net23
rlabel metal1 16422 10778 16422 10778 0 net230
rlabel metal1 19044 14518 19044 14518 0 net231
rlabel metal1 19274 16694 19274 16694 0 net232
rlabel metal1 9890 10166 9890 10166 0 net233
rlabel metal1 10120 22134 10120 22134 0 net234
rlabel metal1 19090 9078 19090 9078 0 net235
rlabel metal2 7590 12517 7590 12517 0 net236
rlabel metal1 19849 10438 19849 10438 0 net237
rlabel metal1 2162 9656 2162 9656 0 net238
rlabel metal1 7682 10234 7682 10234 0 net239
rlabel metal1 13800 2414 13800 2414 0 net24
rlabel metal1 12732 20910 12732 20910 0 net240
rlabel metal2 22908 14212 22908 14212 0 net241
rlabel metal1 23184 4114 23184 4114 0 net242
rlabel metal1 13482 19822 13482 19822 0 net243
rlabel metal1 22816 4794 22816 4794 0 net244
rlabel metal2 21758 6290 21758 6290 0 net245
rlabel metal1 15977 7786 15977 7786 0 net246
rlabel metal2 21206 14042 21206 14042 0 net247
rlabel metal1 22412 15470 22412 15470 0 net248
rlabel metal1 4216 6698 4216 6698 0 net249
rlabel metal1 17388 2414 17388 2414 0 net25
rlabel metal1 16284 5134 16284 5134 0 net250
rlabel metal1 10350 12206 10350 12206 0 net251
rlabel metal1 14025 17170 14025 17170 0 net252
rlabel metal2 18170 13294 18170 13294 0 net253
rlabel metal2 18170 6052 18170 6052 0 net254
rlabel metal1 17112 14042 17112 14042 0 net255
rlabel metal2 16514 14416 16514 14416 0 net256
rlabel metal1 7544 4590 7544 4590 0 net257
rlabel metal1 3726 9554 3726 9554 0 net258
rlabel metal1 2461 9962 2461 9962 0 net259
rlabel metal2 18262 2587 18262 2587 0 net26
rlabel via1 5837 13226 5837 13226 0 net260
rlabel metal1 14158 14382 14158 14382 0 net261
rlabel metal1 7222 4590 7222 4590 0 net262
rlabel metal1 7028 18734 7028 18734 0 net263
rlabel metal1 18538 9078 18538 9078 0 net264
rlabel metal2 22586 14824 22586 14824 0 net265
rlabel metal1 3220 7446 3220 7446 0 net266
rlabel metal1 14137 9622 14137 9622 0 net267
rlabel metal1 3174 14314 3174 14314 0 net268
rlabel metal1 21850 11730 21850 11730 0 net269
rlabel metal1 13018 2448 13018 2448 0 net27
rlabel metal2 17434 5474 17434 5474 0 net270
rlabel metal1 18415 18666 18415 18666 0 net271
rlabel metal1 7033 19346 7033 19346 0 net272
rlabel metal2 19550 6256 19550 6256 0 net273
rlabel metal2 21022 6120 21022 6120 0 net274
rlabel metal1 12844 4590 12844 4590 0 net275
rlabel metal1 5658 7752 5658 7752 0 net276
rlabel metal1 18982 20502 18982 20502 0 net277
rlabel via1 13493 15062 13493 15062 0 net278
rlabel metal1 16095 20910 16095 20910 0 net279
rlabel metal1 6302 2414 6302 2414 0 net28
rlabel metal2 10810 14246 10810 14246 0 net280
rlabel via1 19545 19822 19545 19822 0 net281
rlabel metal1 3772 10166 3772 10166 0 net282
rlabel viali 13482 16558 13482 16558 0 net283
rlabel metal2 3634 14654 3634 14654 0 net284
rlabel metal1 14991 20434 14991 20434 0 net285
rlabel metal1 11316 4114 11316 4114 0 net286
rlabel metal1 5060 17646 5060 17646 0 net287
rlabel metal2 21942 10302 21942 10302 0 net288
rlabel metal1 15773 19414 15773 19414 0 net289
rlabel metal1 7958 2482 7958 2482 0 net29
rlabel metal2 21206 16966 21206 16966 0 net290
rlabel metal1 5504 15402 5504 15402 0 net291
rlabel metal2 4738 17544 4738 17544 0 net292
rlabel metal1 4236 16082 4236 16082 0 net293
rlabel metal2 5106 9350 5106 9350 0 net294
rlabel metal1 14724 9962 14724 9962 0 net295
rlabel via1 8413 19346 8413 19346 0 net296
rlabel metal1 9057 20502 9057 20502 0 net297
rlabel metal2 3358 16694 3358 16694 0 net3
rlabel metal1 5106 10778 5106 10778 0 net30
rlabel metal1 9016 3026 9016 3026 0 net31
rlabel metal1 2070 12138 2070 12138 0 net32
rlabel metal1 2415 14382 2415 14382 0 net33
rlabel metal1 6394 5236 6394 5236 0 net34
rlabel metal1 4232 5882 4232 5882 0 net35
rlabel metal1 2622 6630 2622 6630 0 net36
rlabel metal1 6394 6426 6394 6426 0 net37
rlabel metal1 6164 11730 6164 11730 0 net38
rlabel metal1 3450 15640 3450 15640 0 net39
rlabel metal2 1886 16031 1886 16031 0 net4
rlabel metal1 4830 16116 4830 16116 0 net40
rlabel metal2 1702 14688 1702 14688 0 net41
rlabel metal1 8142 16116 8142 16116 0 net42
rlabel metal1 9430 13430 9430 13430 0 net43
rlabel metal1 8786 19890 8786 19890 0 net44
rlabel metal1 8510 20366 8510 20366 0 net45
rlabel metal1 14122 21046 14122 21046 0 net46
rlabel metal1 13018 20502 13018 20502 0 net47
rlabel metal1 10948 15130 10948 15130 0 net48
rlabel metal1 11914 17714 11914 17714 0 net49
rlabel metal1 11224 24174 11224 24174 0 net5
rlabel metal2 19642 18700 19642 18700 0 net50
rlabel metal1 19136 18802 19136 18802 0 net51
rlabel metal1 19550 14994 19550 14994 0 net52
rlabel metal1 15410 14450 15410 14450 0 net53
rlabel metal1 21620 8602 21620 8602 0 net54
rlabel metal2 23230 15470 23230 15470 0 net55
rlabel metal2 21390 8500 21390 8500 0 net56
rlabel metal1 20700 12886 20700 12886 0 net57
rlabel metal2 21390 6052 21390 6052 0 net58
rlabel metal1 23230 7276 23230 7276 0 net59
rlabel metal2 3082 13498 3082 13498 0 net6
rlabel metal1 16698 6426 16698 6426 0 net60
rlabel metal1 18538 5882 18538 5882 0 net61
rlabel metal1 14168 8602 14168 8602 0 net62
rlabel metal1 13616 12614 13616 12614 0 net63
rlabel metal1 6762 4794 6762 4794 0 net64
rlabel metal1 7406 3706 7406 3706 0 net65
rlabel metal1 6716 5338 6716 5338 0 net66
rlabel metal2 6578 5168 6578 5168 0 net67
rlabel metal1 3128 7514 3128 7514 0 net68
rlabel metal1 9844 3570 9844 3570 0 net69
rlabel metal1 9338 24174 9338 24174 0 net7
rlabel metal1 4232 6834 4232 6834 0 net70
rlabel metal1 6118 13294 6118 13294 0 net71
rlabel metal1 5290 15470 5290 15470 0 net72
rlabel metal1 6394 15028 6394 15028 0 net73
rlabel metal1 9844 17714 9844 17714 0 net74
rlabel metal1 9890 14994 9890 14994 0 net75
rlabel metal1 8510 20468 8510 20468 0 net76
rlabel metal1 8142 19380 8142 19380 0 net77
rlabel metal1 15456 20978 15456 20978 0 net78
rlabel metal1 14582 20434 14582 20434 0 net79
rlabel metal1 7728 24174 7728 24174 0 net8
rlabel metal1 13800 14994 13800 14994 0 net80
rlabel metal2 14398 16422 14398 16422 0 net81
rlabel metal1 18308 18802 18308 18802 0 net82
rlabel metal1 14398 18938 14398 18938 0 net83
rlabel metal1 21022 13906 21022 13906 0 net84
rlabel metal1 18078 14994 18078 14994 0 net85
rlabel metal2 23000 10642 23000 10642 0 net86
rlabel metal1 22954 15538 22954 15538 0 net87
rlabel metal1 21712 5882 21712 5882 0 net88
rlabel metal2 20378 10676 20378 10676 0 net89
rlabel metal1 12788 19958 12788 19958 0 net9
rlabel metal1 23322 5338 23322 5338 0 net90
rlabel metal1 23230 6426 23230 6426 0 net91
rlabel metal1 16192 6426 16192 6426 0 net92
rlabel metal1 16146 7412 16146 7412 0 net93
rlabel metal1 11730 7480 11730 7480 0 net94
rlabel metal1 6210 10234 6210 10234 0 net95
rlabel metal1 7038 4726 7038 4726 0 net96
rlabel metal1 8556 3706 8556 3706 0 net97
rlabel metal1 2208 5338 2208 5338 0 net98
rlabel metal2 3266 7106 3266 7106 0 net99
rlabel metal1 9931 6698 9931 6698 0 regiterFile.memory\[0\]\[0\]
rlabel metal1 3532 14994 3532 14994 0 regiterFile.memory\[0\]\[10\]
rlabel metal1 3532 13906 3532 13906 0 regiterFile.memory\[0\]\[11\]
rlabel metal1 5244 16422 5244 16422 0 regiterFile.memory\[0\]\[12\]
rlabel metal1 6302 13770 6302 13770 0 regiterFile.memory\[0\]\[13\]
rlabel metal1 5198 18938 5198 18938 0 regiterFile.memory\[0\]\[14\]
rlabel metal1 5239 20434 5239 20434 0 regiterFile.memory\[0\]\[15\]
rlabel metal2 10994 21522 10994 21522 0 regiterFile.memory\[0\]\[16\]
rlabel metal2 9614 20196 9614 20196 0 regiterFile.memory\[0\]\[17\]
rlabel metal1 9982 13872 9982 13872 0 regiterFile.memory\[0\]\[18\]
rlabel metal2 12006 17136 12006 17136 0 regiterFile.memory\[0\]\[19\]
rlabel via1 7677 11118 7677 11118 0 regiterFile.memory\[0\]\[1\]
rlabel metal1 16652 17306 16652 17306 0 regiterFile.memory\[0\]\[20\]
rlabel metal1 16560 17850 16560 17850 0 regiterFile.memory\[0\]\[21\]
rlabel metal1 19366 15334 19366 15334 0 regiterFile.memory\[0\]\[22\]
rlabel metal1 14628 12682 14628 12682 0 regiterFile.memory\[0\]\[23\]
rlabel metal1 18211 12818 18211 12818 0 regiterFile.memory\[0\]\[24\]
rlabel metal1 20428 12818 20428 12818 0 regiterFile.memory\[0\]\[25\]
rlabel metal1 19350 9962 19350 9962 0 regiterFile.memory\[0\]\[26\]
rlabel via1 14393 10642 14393 10642 0 regiterFile.memory\[0\]\[27\]
rlabel metal1 18124 7718 18124 7718 0 regiterFile.memory\[0\]\[28\]
rlabel metal1 17705 6698 17705 6698 0 regiterFile.memory\[0\]\[29\]
rlabel metal2 9890 6800 9890 6800 0 regiterFile.memory\[0\]\[2\]
rlabel via1 14393 6766 14393 6766 0 regiterFile.memory\[0\]\[30\]
rlabel metal1 13462 6358 13462 6358 0 regiterFile.memory\[0\]\[31\]
rlabel metal1 10538 4522 10538 4522 0 regiterFile.memory\[0\]\[3\]
rlabel metal1 3082 6256 3082 6256 0 regiterFile.memory\[0\]\[4\]
rlabel metal1 1886 8398 1886 8398 0 regiterFile.memory\[0\]\[5\]
rlabel metal1 4692 7174 4692 7174 0 regiterFile.memory\[0\]\[6\]
rlabel metal1 8678 7446 8678 7446 0 regiterFile.memory\[0\]\[7\]
rlabel via1 3000 12818 3000 12818 0 regiterFile.memory\[0\]\[8\]
rlabel metal1 3496 12410 3496 12410 0 regiterFile.memory\[0\]\[9\]
rlabel metal2 10350 1027 10350 1027 0 rst
<< properties >>
string FIXED_BBOX 0 0 25000 27144
<< end >>
